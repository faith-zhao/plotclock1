module calculate(
	input [7:0] x,
	input [7:0] y,
	output  [31:0] result_1,
	output  [31:0] result_2
);

wire [15:0] xy;
reg [31:0] result1;
reg [31:0] result2;
assign xy = {x[7:0],y[7:0]};
assign result_1 = result1;
assign result_2 = result2;

always@(*) begin
	case(xy)
16'd0 : result1 = 322341;
16'd1 : result1 = 318810;
16'd2 : result1 = 315412;
16'd3 : result1 = 312138;
16'd4 : result1 = 308980;
16'd5 : result1 = 305930;
16'd6 : result1 = 302980;
16'd7 : result1 = 300124;
16'd8 : result1 = 297355;
16'd9 : result1 = 294668;
16'd10 : result1 = 292057;
16'd11 : result1 = 289518;
16'd12 : result1 = 287044;
16'd13 : result1 = 284633;
16'd14 : result1 = 282280;
16'd15 : result1 = 279981;
16'd16 : result1 = 277733;
16'd17 : result1 = 275532;
16'd18 : result1 = 273374;
16'd19 : result1 = 271258;
16'd20 : result1 = 269180;
16'd21 : result1 = 267137;
16'd22 : result1 = 265128;
16'd23 : result1 = 263148;
16'd24 : result1 = 261197;
16'd25 : result1 = 259272;
16'd26 : result1 = 257370;
16'd27 : result1 = 255491;
16'd28 : result1 = 253631;
16'd29 : result1 = 251789;
16'd30 : result1 = 249963;
16'd31 : result1 = 248151;
16'd32 : result1 = 246352;
16'd33 : result1 = 244563;
16'd34 : result1 = 242783;
16'd35 : result1 = 241010;
16'd36 : result1 = 239242;
16'd37 : result1 = 237477;
16'd38 : result1 = 235715;
16'd39 : result1 = 233952;
16'd40 : result1 = 232186;
16'd41 : result1 = 230417;
16'd42 : result1 = 228640;
16'd43 : result1 = 226856;
16'd44 : result1 = 225060;
16'd45 : result1 = 223250;
16'd46 : result1 = 221423;
16'd47 : result1 = 219577;
16'd48 : result1 = 217707;
16'd49 : result1 = 215811;
16'd50 : result1 = 213882;
16'd256 : result1 = 322655;
16'd257 : result1 = 319001;
16'd258 : result1 = 315497;
16'd259 : result1 = 312132;
16'd260 : result1 = 308896;
16'd261 : result1 = 305777;
16'd262 : result1 = 302769;
16'd263 : result1 = 299862;
16'd264 : result1 = 297049;
16'd265 : result1 = 294325;
16'd266 : result1 = 291681;
16'd267 : result1 = 289114;
16'd268 : result1 = 286616;
16'd269 : result1 = 284185;
16'd270 : result1 = 281815;
16'd271 : result1 = 279501;
16'd272 : result1 = 277241;
16'd273 : result1 = 275030;
16'd274 : result1 = 272864;
16'd275 : result1 = 270742;
16'd276 : result1 = 268659;
16'd277 : result1 = 266613;
16'd278 : result1 = 264601;
16'd279 : result1 = 262620;
16'd280 : result1 = 260669;
16'd281 : result1 = 258745;
16'd282 : result1 = 256845;
16'd283 : result1 = 254967;
16'd284 : result1 = 253110;
16'd285 : result1 = 251272;
16'd286 : result1 = 249450;
16'd287 : result1 = 247642;
16'd288 : result1 = 245848;
16'd289 : result1 = 244064;
16'd290 : result1 = 242290;
16'd291 : result1 = 240523;
16'd292 : result1 = 238762;
16'd293 : result1 = 237004;
16'd294 : result1 = 235249;
16'd295 : result1 = 233493;
16'd296 : result1 = 231736;
16'd297 : result1 = 229975;
16'd298 : result1 = 228207;
16'd299 : result1 = 226432;
16'd300 : result1 = 224645;
16'd301 : result1 = 222845;
16'd302 : result1 = 221030;
16'd303 : result1 = 219194;
16'd304 : result1 = 217337;
16'd305 : result1 = 215452;
16'd306 : result1 = 213537;
16'd512 : result1 = 322923;
16'd513 : result1 = 319139;
16'd514 : result1 = 315525;
16'd515 : result1 = 312067;
16'd516 : result1 = 308750;
16'd517 : result1 = 305563;
16'd518 : result1 = 302496;
16'd519 : result1 = 299539;
16'd520 : result1 = 296683;
16'd521 : result1 = 293921;
16'd522 : result1 = 291247;
16'd523 : result1 = 288653;
16'd524 : result1 = 286133;
16'd525 : result1 = 283683;
16'd526 : result1 = 281297;
16'd527 : result1 = 278970;
16'd528 : result1 = 276699;
16'd529 : result1 = 274479;
16'd530 : result1 = 272308;
16'd531 : result1 = 270180;
16'd532 : result1 = 268094;
16'd533 : result1 = 266045;
16'd534 : result1 = 264032;
16'd535 : result1 = 262052;
16'd536 : result1 = 260101;
16'd537 : result1 = 258178;
16'd538 : result1 = 256281;
16'd539 : result1 = 254407;
16'd540 : result1 = 252553;
16'd541 : result1 = 250719;
16'd542 : result1 = 248902;
16'd543 : result1 = 247100;
16'd544 : result1 = 245311;
16'd545 : result1 = 243533;
16'd546 : result1 = 241765;
16'd547 : result1 = 240005;
16'd548 : result1 = 238251;
16'd549 : result1 = 236500;
16'd550 : result1 = 234753;
16'd551 : result1 = 233005;
16'd552 : result1 = 231256;
16'd553 : result1 = 229503;
16'd554 : result1 = 227745;
16'd555 : result1 = 225979;
16'd556 : result1 = 224202;
16'd557 : result1 = 222412;
16'd558 : result1 = 220607;
16'd559 : result1 = 218783;
16'd560 : result1 = 216937;
16'd561 : result1 = 215065;
16'd562 : result1 = 213164;
16'd768 : result1 = 323140;
16'd769 : result1 = 319220;
16'd770 : result1 = 315492;
16'd771 : result1 = 311937;
16'd772 : result1 = 308538;
16'd773 : result1 = 305283;
16'd774 : result1 = 302157;
16'd775 : result1 = 299150;
16'd776 : result1 = 296253;
16'd777 : result1 = 293456;
16'd778 : result1 = 290752;
16'd779 : result1 = 288132;
16'd780 : result1 = 285592;
16'd781 : result1 = 283124;
16'd782 : result1 = 280724;
16'd783 : result1 = 278386;
16'd784 : result1 = 276106;
16'd785 : result1 = 273880;
16'd786 : result1 = 271703;
16'd787 : result1 = 269572;
16'd788 : result1 = 267483;
16'd789 : result1 = 265434;
16'd790 : result1 = 263421;
16'd791 : result1 = 261442;
16'd792 : result1 = 259493;
16'd793 : result1 = 257573;
16'd794 : result1 = 255679;
16'd795 : result1 = 253809;
16'd796 : result1 = 251960;
16'd797 : result1 = 250131;
16'd798 : result1 = 248319;
16'd799 : result1 = 246523;
16'd800 : result1 = 244740;
16'd801 : result1 = 242969;
16'd802 : result1 = 241208;
16'd803 : result1 = 239455;
16'd804 : result1 = 237709;
16'd805 : result1 = 235966;
16'd806 : result1 = 234226;
16'd807 : result1 = 232487;
16'd808 : result1 = 230747;
16'd809 : result1 = 229003;
16'd810 : result1 = 227254;
16'd811 : result1 = 225497;
16'd812 : result1 = 223730;
16'd813 : result1 = 221951;
16'd814 : result1 = 220156;
16'd815 : result1 = 218344;
16'd816 : result1 = 216509;
16'd817 : result1 = 214650;
16'd818 : result1 = 212761;
16'd1024 : result1 = 323300;
16'd1025 : result1 = 319237;
16'd1026 : result1 = 315390;
16'd1027 : result1 = 311737;
16'd1028 : result1 = 308256;
16'd1029 : result1 = 304932;
16'd1030 : result1 = 301749;
16'd1031 : result1 = 298694;
16'd1032 : result1 = 295756;
16'd1033 : result1 = 292926;
16'd1034 : result1 = 290193;
16'd1035 : result1 = 287551;
16'd1036 : result1 = 284992;
16'd1037 : result1 = 282509;
16'd1038 : result1 = 280096;
16'd1039 : result1 = 277749;
16'd1040 : result1 = 275462;
16'd1041 : result1 = 273230;
16'd1042 : result1 = 271049;
16'd1043 : result1 = 268916;
16'd1044 : result1 = 266827;
16'd1045 : result1 = 264778;
16'd1046 : result1 = 262767;
16'd1047 : result1 = 260790;
16'd1048 : result1 = 258845;
16'd1049 : result1 = 256929;
16'd1050 : result1 = 255039;
16'd1051 : result1 = 253174;
16'd1052 : result1 = 251331;
16'd1053 : result1 = 249507;
16'd1054 : result1 = 247702;
16'd1055 : result1 = 245912;
16'd1056 : result1 = 244137;
16'd1057 : result1 = 242373;
16'd1058 : result1 = 240620;
16'd1059 : result1 = 238874;
16'd1060 : result1 = 237136;
16'd1061 : result1 = 235402;
16'd1062 : result1 = 233670;
16'd1063 : result1 = 231940;
16'd1064 : result1 = 230208;
16'd1065 : result1 = 228474;
16'd1066 : result1 = 226734;
16'd1067 : result1 = 224987;
16'd1068 : result1 = 223230;
16'd1069 : result1 = 221461;
16'd1070 : result1 = 219678;
16'd1071 : result1 = 217876;
16'd1072 : result1 = 216053;
16'd1073 : result1 = 214206;
16'd1074 : result1 = 212330;
16'd1280 : result1 = 323396;
16'd1281 : result1 = 319183;
16'd1282 : result1 = 315214;
16'd1283 : result1 = 311461;
16'd1284 : result1 = 307898;
16'd1285 : result1 = 304506;
16'd1286 : result1 = 301266;
16'd1287 : result1 = 298165;
16'd1288 : result1 = 295189;
16'd1289 : result1 = 292327;
16'd1290 : result1 = 289569;
16'd1291 : result1 = 286906;
16'd1292 : result1 = 284330;
16'd1293 : result1 = 281834;
16'd1294 : result1 = 279411;
16'd1295 : result1 = 277056;
16'd1296 : result1 = 274764;
16'd1297 : result1 = 272529;
16'd1298 : result1 = 270346;
16'd1299 : result1 = 268213;
16'd1300 : result1 = 266125;
16'd1301 : result1 = 264078;
16'd1302 : result1 = 262070;
16'd1303 : result1 = 260096;
16'd1304 : result1 = 258156;
16'd1305 : result1 = 256245;
16'd1306 : result1 = 254361;
16'd1307 : result1 = 252501;
16'd1308 : result1 = 250665;
16'd1309 : result1 = 248848;
16'd1310 : result1 = 247050;
16'd1311 : result1 = 245268;
16'd1312 : result1 = 243500;
16'd1313 : result1 = 241744;
16'd1314 : result1 = 239999;
16'd1315 : result1 = 238262;
16'd1316 : result1 = 236532;
16'd1317 : result1 = 234807;
16'd1318 : result1 = 233085;
16'd1319 : result1 = 231363;
16'd1320 : result1 = 229641;
16'd1321 : result1 = 227916;
16'd1322 : result1 = 226186;
16'd1323 : result1 = 224449;
16'd1324 : result1 = 222703;
16'd1325 : result1 = 220944;
16'd1326 : result1 = 219171;
16'd1327 : result1 = 217381;
16'd1328 : result1 = 215570;
16'd1329 : result1 = 213734;
16'd1330 : result1 = 211871;
16'd1536 : result1 = 323420;
16'd1537 : result1 = 319051;
16'd1538 : result1 = 314958;
16'd1539 : result1 = 311103;
16'd1540 : result1 = 307459;
16'd1541 : result1 = 304000;
16'd1542 : result1 = 300706;
16'd1543 : result1 = 297561;
16'd1544 : result1 = 294549;
16'd1545 : result1 = 291658;
16'd1546 : result1 = 288877;
16'd1547 : result1 = 286196;
16'd1548 : result1 = 283606;
16'd1549 : result1 = 281099;
16'd1550 : result1 = 278668;
16'd1551 : result1 = 276308;
16'd1552 : result1 = 274012;
16'd1553 : result1 = 271775;
16'd1554 : result1 = 269593;
16'd1555 : result1 = 267461;
16'd1556 : result1 = 265376;
16'd1557 : result1 = 263333;
16'd1558 : result1 = 261329;
16'd1559 : result1 = 259361;
16'd1560 : result1 = 257425;
16'd1561 : result1 = 255521;
16'd1562 : result1 = 253644;
16'd1563 : result1 = 251792;
16'd1564 : result1 = 249962;
16'd1565 : result1 = 248154;
16'd1566 : result1 = 246364;
16'd1567 : result1 = 244590;
16'd1568 : result1 = 242830;
16'd1569 : result1 = 241083;
16'd1570 : result1 = 239347;
16'd1571 : result1 = 237619;
16'd1572 : result1 = 235898;
16'd1573 : result1 = 234182;
16'd1574 : result1 = 232469;
16'd1575 : result1 = 230758;
16'd1576 : result1 = 229045;
16'd1577 : result1 = 227330;
16'd1578 : result1 = 225610;
16'd1579 : result1 = 223883;
16'd1580 : result1 = 222147;
16'd1581 : result1 = 220399;
16'd1582 : result1 = 218637;
16'd1583 : result1 = 216858;
16'd1584 : result1 = 215058;
16'd1585 : result1 = 213235;
16'd1586 : result1 = 211384;
16'd1792 : result1 = 323364;
16'd1793 : result1 = 318833;
16'd1794 : result1 = 314612;
16'd1795 : result1 = 310657;
16'd1796 : result1 = 306932;
16'd1797 : result1 = 303409;
16'd1798 : result1 = 300064;
16'd1799 : result1 = 296877;
16'd1800 : result1 = 293833;
16'd1801 : result1 = 290916;
16'd1802 : result1 = 288115;
16'd1803 : result1 = 285418;
16'd1804 : result1 = 282816;
16'd1805 : result1 = 280301;
16'd1806 : result1 = 277866;
16'd1807 : result1 = 275502;
16'd1808 : result1 = 273205;
16'd1809 : result1 = 270970;
16'd1810 : result1 = 268790;
16'd1811 : result1 = 266661;
16'd1812 : result1 = 264580;
16'd1813 : result1 = 262542;
16'd1814 : result1 = 260544;
16'd1815 : result1 = 258582;
16'd1816 : result1 = 256654;
16'd1817 : result1 = 254757;
16'd1818 : result1 = 252888;
16'd1819 : result1 = 251044;
16'd1820 : result1 = 249223;
16'd1821 : result1 = 247424;
16'd1822 : result1 = 245642;
16'd1823 : result1 = 243878;
16'd1824 : result1 = 242128;
16'd1825 : result1 = 240390;
16'd1826 : result1 = 238663;
16'd1827 : result1 = 236945;
16'd1828 : result1 = 235234;
16'd1829 : result1 = 233528;
16'd1830 : result1 = 231825;
16'd1831 : result1 = 230123;
16'd1832 : result1 = 228421;
16'd1833 : result1 = 226716;
16'd1834 : result1 = 225006;
16'd1835 : result1 = 223290;
16'd1836 : result1 = 221564;
16'd1837 : result1 = 219827;
16'd1838 : result1 = 218076;
16'd1839 : result1 = 216308;
16'd1840 : result1 = 214520;
16'd1841 : result1 = 212709;
16'd1842 : result1 = 210870;
16'd2048 : result1 = 323218;
16'd2049 : result1 = 318519;
16'd2050 : result1 = 314170;
16'd2051 : result1 = 310115;
16'd2052 : result1 = 306312;
16'd2053 : result1 = 302727;
16'd2054 : result1 = 299334;
16'd2055 : result1 = 296110;
16'd2056 : result1 = 293037;
16'd2057 : result1 = 290098;
16'd2058 : result1 = 287280;
16'd2059 : result1 = 284571;
16'd2060 : result1 = 281961;
16'd2061 : result1 = 279441;
16'd2062 : result1 = 277003;
16'd2063 : result1 = 274639;
16'd2064 : result1 = 272343;
16'd2065 : result1 = 270110;
16'd2066 : result1 = 267935;
16'd2067 : result1 = 265811;
16'd2068 : result1 = 263736;
16'd2069 : result1 = 261705;
16'd2070 : result1 = 259715;
16'd2071 : result1 = 257761;
16'd2072 : result1 = 255842;
16'd2073 : result1 = 253954;
16'd2074 : result1 = 252093;
16'd2075 : result1 = 250259;
16'd2076 : result1 = 248448;
16'd2077 : result1 = 246658;
16'd2078 : result1 = 244887;
16'd2079 : result1 = 243132;
16'd2080 : result1 = 241392;
16'd2081 : result1 = 239665;
16'd2082 : result1 = 237948;
16'd2083 : result1 = 236240;
16'd2084 : result1 = 234539;
16'd2085 : result1 = 232844;
16'd2086 : result1 = 231151;
16'd2087 : result1 = 229460;
16'd2088 : result1 = 227768;
16'd2089 : result1 = 226074;
16'd2090 : result1 = 224375;
16'd2091 : result1 = 222669;
16'd2092 : result1 = 220954;
16'd2093 : result1 = 219228;
16'd2094 : result1 = 217488;
16'd2095 : result1 = 215732;
16'd2096 : result1 = 213955;
16'd2097 : result1 = 212156;
16'd2098 : result1 = 210329;
16'd2304 : result1 = 322968;
16'd2305 : result1 = 318099;
16'd2306 : result1 = 313622;
16'd2307 : result1 = 309470;
16'd2308 : result1 = 305593;
16'd2309 : result1 = 301951;
16'd2310 : result1 = 298514;
16'd2311 : result1 = 295257;
16'd2312 : result1 = 292158;
16'd2313 : result1 = 289201;
16'd2314 : result1 = 286370;
16'd2315 : result1 = 283653;
16'd2316 : result1 = 281038;
16'd2317 : result1 = 278516;
16'd2318 : result1 = 276078;
16'd2319 : result1 = 273717;
16'd2320 : result1 = 271425;
16'd2321 : result1 = 269197;
16'd2322 : result1 = 267028;
16'd2323 : result1 = 264912;
16'd2324 : result1 = 262845;
16'd2325 : result1 = 260823;
16'd2326 : result1 = 258842;
16'd2327 : result1 = 256898;
16'd2328 : result1 = 254988;
16'd2329 : result1 = 253110;
16'd2330 : result1 = 251261;
16'd2331 : result1 = 249437;
16'd2332 : result1 = 247637;
16'd2333 : result1 = 245857;
16'd2334 : result1 = 244097;
16'd2335 : result1 = 242353;
16'd2336 : result1 = 240624;
16'd2337 : result1 = 238908;
16'd2338 : result1 = 237202;
16'd2339 : result1 = 235505;
16'd2340 : result1 = 233815;
16'd2341 : result1 = 232130;
16'd2342 : result1 = 230448;
16'd2343 : result1 = 228768;
16'd2344 : result1 = 227087;
16'd2345 : result1 = 225404;
16'd2346 : result1 = 223716;
16'd2347 : result1 = 222021;
16'd2348 : result1 = 220318;
16'd2349 : result1 = 218603;
16'd2350 : result1 = 216874;
16'd2351 : result1 = 215129;
16'd2352 : result1 = 213364;
16'd2353 : result1 = 211576;
16'd2354 : result1 = 209762;
16'd2560 : result1 = 322603;
16'd2561 : result1 = 317562;
16'd2562 : result1 = 312959;
16'd2563 : result1 = 308714;
16'd2564 : result1 = 304767;
16'd2565 : result1 = 301074;
16'd2566 : result1 = 297599;
16'd2567 : result1 = 294313;
16'd2568 : result1 = 291195;
16'd2569 : result1 = 288224;
16'd2570 : result1 = 285384;
16'd2571 : result1 = 282662;
16'd2572 : result1 = 280046;
16'd2573 : result1 = 277525;
16'd2574 : result1 = 275091;
16'd2575 : result1 = 272735;
16'd2576 : result1 = 270450;
16'd2577 : result1 = 268230;
16'd2578 : result1 = 266070;
16'd2579 : result1 = 263963;
16'd2580 : result1 = 261906;
16'd2581 : result1 = 259895;
16'd2582 : result1 = 257924;
16'd2583 : result1 = 255992;
16'd2584 : result1 = 254094;
16'd2585 : result1 = 252227;
16'd2586 : result1 = 250389;
16'd2587 : result1 = 248577;
16'd2588 : result1 = 246789;
16'd2589 : result1 = 245021;
16'd2590 : result1 = 243273;
16'd2591 : result1 = 241541;
16'd2592 : result1 = 239824;
16'd2593 : result1 = 238119;
16'd2594 : result1 = 236425;
16'd2595 : result1 = 234739;
16'd2596 : result1 = 233061;
16'd2597 : result1 = 231388;
16'd2598 : result1 = 229717;
16'd2599 : result1 = 228048;
16'd2600 : result1 = 226379;
16'd2601 : result1 = 224707;
16'd2602 : result1 = 223030;
16'd2603 : result1 = 221346;
16'd2604 : result1 = 219654;
16'd2605 : result1 = 217951;
16'd2606 : result1 = 216233;
16'd2607 : result1 = 214500;
16'd2608 : result1 = 212747;
16'd2609 : result1 = 210971;
16'd2610 : result1 = 209168;
16'd2816 : result1 = 322108;
16'd2817 : result1 = 316895;
16'd2818 : result1 = 312172;
16'd2819 : result1 = 307840;
16'd2820 : result1 = 303830;
16'd2821 : result1 = 300092;
16'd2822 : result1 = 296584;
16'd2823 : result1 = 293276;
16'd2824 : result1 = 290143;
16'd2825 : result1 = 287164;
16'd2826 : result1 = 284320;
16'd2827 : result1 = 281598;
16'd2828 : result1 = 278984;
16'd2829 : result1 = 276469;
16'd2830 : result1 = 274041;
16'd2831 : result1 = 271693;
16'd2832 : result1 = 269418;
16'd2833 : result1 = 267209;
16'd2834 : result1 = 265059;
16'd2835 : result1 = 262965;
16'd2836 : result1 = 260920;
16'd2837 : result1 = 258921;
16'd2838 : result1 = 256963;
16'd2839 : result1 = 255043;
16'd2840 : result1 = 253158;
16'd2841 : result1 = 251305;
16'd2842 : result1 = 249480;
16'd2843 : result1 = 247681;
16'd2844 : result1 = 245905;
16'd2845 : result1 = 244151;
16'd2846 : result1 = 242415;
16'd2847 : result1 = 240696;
16'd2848 : result1 = 238991;
16'd2849 : result1 = 237299;
16'd2850 : result1 = 235617;
16'd2851 : result1 = 233944;
16'd2852 : result1 = 232277;
16'd2853 : result1 = 230616;
16'd2854 : result1 = 228958;
16'd2855 : result1 = 227301;
16'd2856 : result1 = 225643;
16'd2857 : result1 = 223982;
16'd2858 : result1 = 222317;
16'd2859 : result1 = 220645;
16'd2860 : result1 = 218965;
16'd2861 : result1 = 217273;
16'd2862 : result1 = 215567;
16'd2863 : result1 = 213845;
16'd2864 : result1 = 212103;
16'd2865 : result1 = 210339;
16'd2866 : result1 = 208549;
16'd3072 : result1 = 321465;
16'd3073 : result1 = 316087;
16'd3074 : result1 = 311250;
16'd3075 : result1 = 306840;
16'd3076 : result1 = 302775;
16'd3077 : result1 = 298999;
16'd3078 : result1 = 295467;
16'd3079 : result1 = 292143;
16'd3080 : result1 = 289002;
16'd3081 : result1 = 286019;
16'd3082 : result1 = 283176;
16'd3083 : result1 = 280458;
16'd3084 : result1 = 277852;
16'd3085 : result1 = 275345;
16'd3086 : result1 = 272928;
16'd3087 : result1 = 270592;
16'd3088 : result1 = 268329;
16'd3089 : result1 = 266133;
16'd3090 : result1 = 263997;
16'd3091 : result1 = 261916;
16'd3092 : result1 = 259886;
16'd3093 : result1 = 257901;
16'd3094 : result1 = 255958;
16'd3095 : result1 = 254053;
16'd3096 : result1 = 252182;
16'd3097 : result1 = 250343;
16'd3098 : result1 = 248533;
16'd3099 : result1 = 246748;
16'd3100 : result1 = 244986;
16'd3101 : result1 = 243246;
16'd3102 : result1 = 241523;
16'd3103 : result1 = 239818;
16'd3104 : result1 = 238126;
16'd3105 : result1 = 236447;
16'd3106 : result1 = 234779;
16'd3107 : result1 = 233118;
16'd3108 : result1 = 231465;
16'd3109 : result1 = 229816;
16'd3110 : result1 = 228170;
16'd3111 : result1 = 226525;
16'd3112 : result1 = 224880;
16'd3113 : result1 = 223231;
16'd3114 : result1 = 221578;
16'd3115 : result1 = 219918;
16'd3116 : result1 = 218249;
16'd3117 : result1 = 216569;
16'd3118 : result1 = 214875;
16'd3119 : result1 = 213164;
16'd3120 : result1 = 211435;
16'd3121 : result1 = 209682;
16'd3122 : result1 = 207904;
16'd3328 : result1 = 320659;
16'd3329 : result1 = 315123;
16'd3330 : result1 = 310184;
16'd3331 : result1 = 305706;
16'd3332 : result1 = 301597;
16'd3333 : result1 = 297792;
16'd3334 : result1 = 294243;
16'd3335 : result1 = 290911;
16'd3336 : result1 = 287768;
16'd3337 : result1 = 284788;
16'd3338 : result1 = 281952;
16'd3339 : result1 = 279244;
16'd3340 : result1 = 276648;
16'd3341 : result1 = 274154;
16'd3342 : result1 = 271751;
16'd3343 : result1 = 269430;
16'd3344 : result1 = 267183;
16'd3345 : result1 = 265002;
16'd3346 : result1 = 262883;
16'd3347 : result1 = 260818;
16'd3348 : result1 = 258804;
16'd3349 : result1 = 256836;
16'd3350 : result1 = 254909;
16'd3351 : result1 = 253020;
16'd3352 : result1 = 251166;
16'd3353 : result1 = 249342;
16'd3354 : result1 = 247548;
16'd3355 : result1 = 245778;
16'd3356 : result1 = 244032;
16'd3357 : result1 = 242306;
16'd3358 : result1 = 240599;
16'd3359 : result1 = 238908;
16'd3360 : result1 = 237230;
16'd3361 : result1 = 235565;
16'd3362 : result1 = 233910;
16'd3363 : result1 = 232264;
16'd3364 : result1 = 230623;
16'd3365 : result1 = 228988;
16'd3366 : result1 = 227355;
16'd3367 : result1 = 225723;
16'd3368 : result1 = 224090;
16'd3369 : result1 = 222454;
16'd3370 : result1 = 220813;
16'd3371 : result1 = 219165;
16'd3372 : result1 = 217508;
16'd3373 : result1 = 215839;
16'd3374 : result1 = 214157;
16'd3375 : result1 = 212459;
16'd3376 : result1 = 210741;
16'd3377 : result1 = 209001;
16'd3378 : result1 = 207234;
16'd3584 : result1 = 319669;
16'd3585 : result1 = 313991;
16'd3586 : result1 = 308964;
16'd3587 : result1 = 304431;
16'd3588 : result1 = 300289;
16'd3589 : result1 = 296467;
16'd3590 : result1 = 292910;
16'd3591 : result1 = 289579;
16'd3592 : result1 = 286441;
16'd3593 : result1 = 283470;
16'd3594 : result1 = 280647;
16'd3595 : result1 = 277952;
16'd3596 : result1 = 275373;
16'd3597 : result1 = 272896;
16'd3598 : result1 = 270511;
16'd3599 : result1 = 268208;
16'd3600 : result1 = 265979;
16'd3601 : result1 = 263818;
16'd3602 : result1 = 261717;
16'd3603 : result1 = 259671;
16'd3604 : result1 = 257676;
16'd3605 : result1 = 255726;
16'd3606 : result1 = 253817;
16'd3607 : result1 = 251946;
16'd3608 : result1 = 250109;
16'd3609 : result1 = 248303;
16'd3610 : result1 = 246525;
16'd3611 : result1 = 244773;
16'd3612 : result1 = 243043;
16'd3613 : result1 = 241333;
16'd3614 : result1 = 239641;
16'd3615 : result1 = 237965;
16'd3616 : result1 = 236303;
16'd3617 : result1 = 234653;
16'd3618 : result1 = 233013;
16'd3619 : result1 = 231380;
16'd3620 : result1 = 229754;
16'd3621 : result1 = 228132;
16'd3622 : result1 = 226512;
16'd3623 : result1 = 224893;
16'd3624 : result1 = 223273;
16'd3625 : result1 = 221650;
16'd3626 : result1 = 220021;
16'd3627 : result1 = 218386;
16'd3628 : result1 = 216741;
16'd3629 : result1 = 215085;
16'd3630 : result1 = 213415;
16'd3631 : result1 = 211728;
16'd3632 : result1 = 210022;
16'd3633 : result1 = 208294;
16'd3634 : result1 = 206539;
16'd3840 : result1 = 318478;
16'd3841 : result1 = 312678;
16'd3842 : result1 = 307581;
16'd3843 : result1 = 303010;
16'd3844 : result1 = 298849;
16'd3845 : result1 = 295020;
16'd3846 : result1 = 291466;
16'd3847 : result1 = 288144;
16'd3848 : result1 = 285019;
16'd3849 : result1 = 282065;
16'd3850 : result1 = 279260;
16'd3851 : result1 = 276585;
16'd3852 : result1 = 274027;
16'd3853 : result1 = 271571;
16'd3854 : result1 = 269208;
16'd3855 : result1 = 266927;
16'd3856 : result1 = 264720;
16'd3857 : result1 = 262580;
16'd3858 : result1 = 260500;
16'd3859 : result1 = 258476;
16'd3860 : result1 = 256501;
16'd3861 : result1 = 254572;
16'd3862 : result1 = 252683;
16'd3863 : result1 = 250831;
16'd3864 : result1 = 249014;
16'd3865 : result1 = 247226;
16'd3866 : result1 = 245467;
16'd3867 : result1 = 243732;
16'd3868 : result1 = 242019;
16'd3869 : result1 = 240327;
16'd3870 : result1 = 238651;
16'd3871 : result1 = 236992;
16'd3872 : result1 = 235346;
16'd3873 : result1 = 233711;
16'd3874 : result1 = 232086;
16'd3875 : result1 = 230468;
16'd3876 : result1 = 228856;
16'd3877 : result1 = 227248;
16'd3878 : result1 = 225642;
16'd3879 : result1 = 224037;
16'd3880 : result1 = 222430;
16'd3881 : result1 = 220820;
16'd3882 : result1 = 219205;
16'd3883 : result1 = 217582;
16'd3884 : result1 = 215950;
16'd3885 : result1 = 214306;
16'd3886 : result1 = 212648;
16'd3887 : result1 = 210973;
16'd3888 : result1 = 209279;
16'd3889 : result1 = 207563;
16'd3890 : result1 = 205820;
16'd4096 : result1 = 317066;
16'd4097 : result1 = 311172;
16'd4098 : result1 = 306028;
16'd4099 : result1 = 301436;
16'd4100 : result1 = 297272;
16'd4101 : result1 = 293450;
16'd4102 : result1 = 289910;
16'd4103 : result1 = 286606;
16'd4104 : result1 = 283503;
16'd4105 : result1 = 280572;
16'd4106 : result1 = 277791;
16'd4107 : result1 = 275142;
16'd4108 : result1 = 272610;
16'd4109 : result1 = 270180;
16'd4110 : result1 = 267842;
16'd4111 : result1 = 265586;
16'd4112 : result1 = 263404;
16'd4113 : result1 = 261289;
16'd4114 : result1 = 259234;
16'd4115 : result1 = 257233;
16'd4116 : result1 = 255281;
16'd4117 : result1 = 253373;
16'd4118 : result1 = 251507;
16'd4119 : result1 = 249676;
16'd4120 : result1 = 247879;
16'd4121 : result1 = 246112;
16'd4122 : result1 = 244372;
16'd4123 : result1 = 242656;
16'd4124 : result1 = 240962;
16'd4125 : result1 = 239287;
16'd4126 : result1 = 237630;
16'd4127 : result1 = 235987;
16'd4128 : result1 = 234358;
16'd4129 : result1 = 232739;
16'd4130 : result1 = 231130;
16'd4131 : result1 = 229527;
16'd4132 : result1 = 227931;
16'd4133 : result1 = 226338;
16'd4134 : result1 = 224746;
16'd4135 : result1 = 223155;
16'd4136 : result1 = 221562;
16'd4137 : result1 = 219965;
16'd4138 : result1 = 218363;
16'd4139 : result1 = 216753;
16'd4140 : result1 = 215134;
16'd4141 : result1 = 213502;
16'd4142 : result1 = 211857;
16'd4143 : result1 = 210194;
16'd4144 : result1 = 208512;
16'd4145 : result1 = 206807;
16'd4146 : result1 = 205076;
16'd4352 : result1 = 315418;
16'd4353 : result1 = 309463;
16'd4354 : result1 = 304299;
16'd4355 : result1 = 299708;
16'd4356 : result1 = 295557;
16'd4357 : result1 = 291756;
16'd4358 : result1 = 288241;
16'd4359 : result1 = 284965;
16'd4360 : result1 = 281892;
16'd4361 : result1 = 278992;
16'd4362 : result1 = 276242;
16'd4363 : result1 = 273624;
16'd4364 : result1 = 271122;
16'd4365 : result1 = 268723;
16'd4366 : result1 = 266414;
16'd4367 : result1 = 264188;
16'd4368 : result1 = 262034;
16'd4369 : result1 = 259946;
16'd4370 : result1 = 257917;
16'd4371 : result1 = 255942;
16'd4372 : result1 = 254015;
16'd4373 : result1 = 252132;
16'd4374 : result1 = 250289;
16'd4375 : result1 = 248482;
16'd4376 : result1 = 246707;
16'd4377 : result1 = 244961;
16'd4378 : result1 = 243242;
16'd4379 : result1 = 241546;
16'd4380 : result1 = 239872;
16'd4381 : result1 = 238216;
16'd4382 : result1 = 236577;
16'd4383 : result1 = 234952;
16'd4384 : result1 = 233340;
16'd4385 : result1 = 231739;
16'd4386 : result1 = 230146;
16'd4387 : result1 = 228559;
16'd4388 : result1 = 226978;
16'd4389 : result1 = 225400;
16'd4390 : result1 = 223824;
16'd4391 : result1 = 222247;
16'd4392 : result1 = 220668;
16'd4393 : result1 = 219085;
16'd4394 : result1 = 217496;
16'd4395 : result1 = 215900;
16'd4396 : result1 = 214293;
16'd4397 : result1 = 212674;
16'd4398 : result1 = 211041;
16'd4399 : result1 = 209391;
16'd4400 : result1 = 207721;
16'd4401 : result1 = 206028;
16'd4402 : result1 = 204309;
16'd4608 : result1 = 313520;
16'd4609 : result1 = 307546;
16'd4610 : result1 = 302390;
16'd4611 : result1 = 297822;
16'd4612 : result1 = 293702;
16'd4613 : result1 = 289937;
16'd4614 : result1 = 286460;
16'd4615 : result1 = 283222;
16'd4616 : result1 = 280187;
16'd4617 : result1 = 277326;
16'd4618 : result1 = 274614;
16'd4619 : result1 = 272033;
16'd4620 : result1 = 269566;
16'd4621 : result1 = 267201;
16'd4622 : result1 = 264927;
16'd4623 : result1 = 262732;
16'd4624 : result1 = 260610;
16'd4625 : result1 = 258552;
16'd4626 : result1 = 256552;
16'd4627 : result1 = 254605;
16'd4628 : result1 = 252706;
16'd4629 : result1 = 250849;
16'd4630 : result1 = 249031;
16'd4631 : result1 = 247248;
16'd4632 : result1 = 245497;
16'd4633 : result1 = 243774;
16'd4634 : result1 = 242077;
16'd4635 : result1 = 240402;
16'd4636 : result1 = 238749;
16'd4637 : result1 = 237113;
16'd4638 : result1 = 235493;
16'd4639 : result1 = 233887;
16'd4640 : result1 = 232294;
16'd4641 : result1 = 230710;
16'd4642 : result1 = 229134;
16'd4643 : result1 = 227564;
16'd4644 : result1 = 225999;
16'd4645 : result1 = 224437;
16'd4646 : result1 = 222876;
16'd4647 : result1 = 221314;
16'd4648 : result1 = 219749;
16'd4649 : result1 = 218181;
16'd4650 : result1 = 216606;
16'd4651 : result1 = 215022;
16'd4652 : result1 = 213429;
16'd4653 : result1 = 211823;
16'd4654 : result1 = 210202;
16'd4655 : result1 = 208564;
16'd4656 : result1 = 206906;
16'd4657 : result1 = 205225;
16'd4658 : result1 = 203517;
16'd4864 : result1 = 311363;
16'd4865 : result1 = 305415;
16'd4866 : result1 = 300300;
16'd4867 : result1 = 295779;
16'd4868 : result1 = 291709;
16'd4869 : result1 = 287994;
16'd4870 : result1 = 284567;
16'd4871 : result1 = 281379;
16'd4872 : result1 = 278391;
16'd4873 : result1 = 275575;
16'd4874 : result1 = 272908;
16'd4875 : result1 = 270369;
16'd4876 : result1 = 267943;
16'd4877 : result1 = 265617;
16'd4878 : result1 = 263380;
16'd4879 : result1 = 261221;
16'd4880 : result1 = 259133;
16'd4881 : result1 = 257108;
16'd4882 : result1 = 255140;
16'd4883 : result1 = 253224;
16'd4884 : result1 = 251353;
16'd4885 : result1 = 249525;
16'd4886 : result1 = 247734;
16'd4887 : result1 = 245977;
16'd4888 : result1 = 244250;
16'd4889 : result1 = 242552;
16'd4890 : result1 = 240878;
16'd4891 : result1 = 239226;
16'd4892 : result1 = 237594;
16'd4893 : result1 = 235979;
16'd4894 : result1 = 234380;
16'd4895 : result1 = 232793;
16'd4896 : result1 = 231218;
16'd4897 : result1 = 229653;
16'd4898 : result1 = 228095;
16'd4899 : result1 = 226542;
16'd4900 : result1 = 224994;
16'd4901 : result1 = 223448;
16'd4902 : result1 = 221902;
16'd4903 : result1 = 220356;
16'd4904 : result1 = 218806;
16'd4905 : result1 = 217252;
16'd4906 : result1 = 215691;
16'd4907 : result1 = 214121;
16'd4908 : result1 = 212541;
16'd4909 : result1 = 210948;
16'd4910 : result1 = 209340;
16'd4911 : result1 = 207714;
16'd4912 : result1 = 206068;
16'd4913 : result1 = 204399;
16'd4914 : result1 = 202703;
16'd5120 : result1 = 308946;
16'd5121 : result1 = 303072;
16'd5122 : result1 = 298030;
16'd5123 : result1 = 293582;
16'd5124 : result1 = 289581;
16'd5125 : result1 = 285932;
16'd5126 : result1 = 282567;
16'd5127 : result1 = 279437;
16'd5128 : result1 = 276506;
16'd5129 : result1 = 273743;
16'd5130 : result1 = 271126;
16'd5131 : result1 = 268635;
16'd5132 : result1 = 266254;
16'd5133 : result1 = 263972;
16'd5134 : result1 = 261775;
16'd5135 : result1 = 259656;
16'd5136 : result1 = 257605;
16'd5137 : result1 = 255616;
16'd5138 : result1 = 253682;
16'd5139 : result1 = 251798;
16'd5140 : result1 = 249959;
16'd5141 : result1 = 248161;
16'd5142 : result1 = 246398;
16'd5143 : result1 = 244669;
16'd5144 : result1 = 242969;
16'd5145 : result1 = 241295;
16'd5146 : result1 = 239646;
16'd5147 : result1 = 238018;
16'd5148 : result1 = 236408;
16'd5149 : result1 = 234815;
16'd5150 : result1 = 233237;
16'd5151 : result1 = 231671;
16'd5152 : result1 = 230115;
16'd5153 : result1 = 228569;
16'd5154 : result1 = 227029;
16'd5155 : result1 = 225494;
16'd5156 : result1 = 223963;
16'd5157 : result1 = 222434;
16'd5158 : result1 = 220904;
16'd5159 : result1 = 219373;
16'd5160 : result1 = 217839;
16'd5161 : result1 = 216299;
16'd5162 : result1 = 214752;
16'd5163 : result1 = 213197;
16'd5164 : result1 = 211630;
16'd5165 : result1 = 210050;
16'd5166 : result1 = 208455;
16'd5167 : result1 = 206842;
16'd5168 : result1 = 205208;
16'd5169 : result1 = 203550;
16'd5170 : result1 = 201866;
16'd5376 : result1 = 306274;
16'd5377 : result1 = 300521;
16'd5378 : result1 = 295587;
16'd5379 : result1 = 291234;
16'd5380 : result1 = 287321;
16'd5381 : result1 = 283752;
16'd5382 : result1 = 280462;
16'd5383 : result1 = 277402;
16'd5384 : result1 = 274535;
16'd5385 : result1 = 271832;
16'd5386 : result1 = 269271;
16'd5387 : result1 = 266833;
16'd5388 : result1 = 264503;
16'd5389 : result1 = 262268;
16'd5390 : result1 = 260116;
16'd5391 : result1 = 258039;
16'd5392 : result1 = 256028;
16'd5393 : result1 = 254078;
16'd5394 : result1 = 252180;
16'd5395 : result1 = 250331;
16'd5396 : result1 = 248525;
16'd5397 : result1 = 246758;
16'd5398 : result1 = 245025;
16'd5399 : result1 = 243325;
16'd5400 : result1 = 241653;
16'd5401 : result1 = 240006;
16'd5402 : result1 = 238382;
16'd5403 : result1 = 236778;
16'd5404 : result1 = 235192;
16'd5405 : result1 = 233622;
16'd5406 : result1 = 232065;
16'd5407 : result1 = 230520;
16'd5408 : result1 = 228985;
16'd5409 : result1 = 227458;
16'd5410 : result1 = 225937;
16'd5411 : result1 = 224421;
16'd5412 : result1 = 222907;
16'd5413 : result1 = 221395;
16'd5414 : result1 = 219882;
16'd5415 : result1 = 218367;
16'd5416 : result1 = 216848;
16'd5417 : result1 = 215323;
16'd5418 : result1 = 213791;
16'd5419 : result1 = 212249;
16'd5420 : result1 = 210696;
16'd5421 : result1 = 209129;
16'd5422 : result1 = 207547;
16'd5423 : result1 = 205946;
16'd5424 : result1 = 204325;
16'd5425 : result1 = 202679;
16'd5426 : result1 = 201006;
16'd5632 : result1 = 303356;
16'd5633 : result1 = 297772;
16'd5634 : result1 = 292977;
16'd5635 : result1 = 288744;
16'd5636 : result1 = 284936;
16'd5637 : result1 = 281462;
16'd5638 : result1 = 278257;
16'd5639 : result1 = 275276;
16'd5640 : result1 = 272481;
16'd5641 : result1 = 269845;
16'd5642 : result1 = 267347;
16'd5643 : result1 = 264967;
16'd5644 : result1 = 262691;
16'd5645 : result1 = 260507;
16'd5646 : result1 = 258403;
16'd5647 : result1 = 256372;
16'd5648 : result1 = 254404;
16'd5649 : result1 = 252494;
16'd5650 : result1 = 250635;
16'd5651 : result1 = 248823;
16'd5652 : result1 = 247051;
16'd5653 : result1 = 245317;
16'd5654 : result1 = 243617;
16'd5655 : result1 = 241947;
16'd5656 : result1 = 240303;
16'd5657 : result1 = 238684;
16'd5658 : result1 = 237087;
16'd5659 : result1 = 235508;
16'd5660 : result1 = 233947;
16'd5661 : result1 = 232400;
16'd5662 : result1 = 230866;
16'd5663 : result1 = 229343;
16'd5664 : result1 = 227828;
16'd5665 : result1 = 226321;
16'd5666 : result1 = 224820;
16'd5667 : result1 = 223322;
16'd5668 : result1 = 221826;
16'd5669 : result1 = 220332;
16'd5670 : result1 = 218835;
16'd5671 : result1 = 217337;
16'd5672 : result1 = 215833;
16'd5673 : result1 = 214324;
16'd5674 : result1 = 212806;
16'd5675 : result1 = 211279;
16'd5676 : result1 = 209740;
16'd5677 : result1 = 208186;
16'd5678 : result1 = 206617;
16'd5679 : result1 = 205029;
16'd5680 : result1 = 203419;
16'd5681 : result1 = 201785;
16'd5682 : result1 = 200123;
16'd5888 : result1 = 300213;
16'd5889 : result1 = 294838;
16'd5890 : result1 = 290211;
16'd5891 : result1 = 286119;
16'd5892 : result1 = 282433;
16'd5893 : result1 = 279067;
16'd5894 : result1 = 275959;
16'd5895 : result1 = 273065;
16'd5896 : result1 = 270350;
16'd5897 : result1 = 267787;
16'd5898 : result1 = 265357;
16'd5899 : result1 = 263040;
16'd5900 : result1 = 260822;
16'd5901 : result1 = 258693;
16'd5902 : result1 = 256640;
16'd5903 : result1 = 254657;
16'd5904 : result1 = 252735;
16'd5905 : result1 = 250868;
16'd5906 : result1 = 249049;
16'd5907 : result1 = 247275;
16'd5908 : result1 = 245540;
16'd5909 : result1 = 243841;
16'd5910 : result1 = 242174;
16'd5911 : result1 = 240535;
16'd5912 : result1 = 238922;
16'd5913 : result1 = 237331;
16'd5914 : result1 = 235761;
16'd5915 : result1 = 234209;
16'd5916 : result1 = 232673;
16'd5917 : result1 = 231150;
16'd5918 : result1 = 229640;
16'd5919 : result1 = 228139;
16'd5920 : result1 = 226646;
16'd5921 : result1 = 225159;
16'd5922 : result1 = 223678;
16'd5923 : result1 = 222199;
16'd5924 : result1 = 220722;
16'd5925 : result1 = 219245;
16'd5926 : result1 = 217766;
16'd5927 : result1 = 216284;
16'd5928 : result1 = 214796;
16'd5929 : result1 = 213302;
16'd5930 : result1 = 211800;
16'd5931 : result1 = 210287;
16'd5932 : result1 = 208761;
16'd5933 : result1 = 207222;
16'd5934 : result1 = 205665;
16'd5935 : result1 = 204089;
16'd5936 : result1 = 202492;
16'd5937 : result1 = 200869;
16'd5938 : result1 = 199219;
16'd6144 : result1 = 296867;
16'd6145 : result1 = 291738;
16'd6146 : result1 = 287303;
16'd6147 : result1 = 283371;
16'd6148 : result1 = 279822;
16'd6149 : result1 = 276575;
16'd6150 : result1 = 273573;
16'd6151 : result1 = 270774;
16'd6152 : result1 = 268146;
16'd6153 : result1 = 265663;
16'd6154 : result1 = 263304;
16'd6155 : result1 = 261054;
16'd6156 : result1 = 258899;
16'd6157 : result1 = 256828;
16'd6158 : result1 = 254830;
16'd6159 : result1 = 252897;
16'd6160 : result1 = 251023;
16'd6161 : result1 = 249200;
16'd6162 : result1 = 247425;
16'd6163 : result1 = 245691;
16'd6164 : result1 = 243994;
16'd6165 : result1 = 242331;
16'd6166 : result1 = 240698;
16'd6167 : result1 = 239092;
16'd6168 : result1 = 237509;
16'd6169 : result1 = 235949;
16'd6170 : result1 = 234407;
16'd6171 : result1 = 232882;
16'd6172 : result1 = 231372;
16'd6173 : result1 = 229874;
16'd6174 : result1 = 228387;
16'd6175 : result1 = 226909;
16'd6176 : result1 = 225438;
16'd6177 : result1 = 223973;
16'd6178 : result1 = 222512;
16'd6179 : result1 = 221053;
16'd6180 : result1 = 219594;
16'd6181 : result1 = 218135;
16'd6182 : result1 = 216674;
16'd6183 : result1 = 215208;
16'd6184 : result1 = 213737;
16'd6185 : result1 = 212259;
16'd6186 : result1 = 210771;
16'd6187 : result1 = 209273;
16'd6188 : result1 = 207762;
16'd6189 : result1 = 206235;
16'd6190 : result1 = 204692;
16'd6191 : result1 = 203129;
16'd6192 : result1 = 201543;
16'd6193 : result1 = 199932;
16'd6194 : result1 = 198293;
16'd6400 : result1 = 293347;
16'd6401 : result1 = 288490;
16'd6402 : result1 = 284269;
16'd6403 : result1 = 280513;
16'd6404 : result1 = 277113;
16'd6405 : result1 = 273995;
16'd6406 : result1 = 271108;
16'd6407 : result1 = 268411;
16'd6408 : result1 = 265875;
16'd6409 : result1 = 263476;
16'd6410 : result1 = 261195;
16'd6411 : result1 = 259016;
16'd6412 : result1 = 256926;
16'd6413 : result1 = 254915;
16'd6414 : result1 = 252974;
16'd6415 : result1 = 251095;
16'd6416 : result1 = 249270;
16'd6417 : result1 = 247495;
16'd6418 : result1 = 245763;
16'd6419 : result1 = 244071;
16'd6420 : result1 = 242413;
16'd6421 : result1 = 240788;
16'd6422 : result1 = 239190;
16'd6423 : result1 = 237618;
16'd6424 : result1 = 236068;
16'd6425 : result1 = 234537;
16'd6426 : result1 = 233025;
16'd6427 : result1 = 231528;
16'd6428 : result1 = 230044;
16'd6429 : result1 = 228572;
16'd6430 : result1 = 227109;
16'd6431 : result1 = 225655;
16'd6432 : result1 = 224206;
16'd6433 : result1 = 222763;
16'd6434 : result1 = 221322;
16'd6435 : result1 = 219883;
16'd6436 : result1 = 218444;
16'd6437 : result1 = 217003;
16'd6438 : result1 = 215560;
16'd6439 : result1 = 214111;
16'd6440 : result1 = 212656;
16'd6441 : result1 = 211194;
16'd6442 : result1 = 209721;
16'd6443 : result1 = 208238;
16'd6444 : result1 = 206740;
16'd6445 : result1 = 205228;
16'd6446 : result1 = 203697;
16'd6447 : result1 = 202146;
16'd6448 : result1 = 200573;
16'd6449 : result1 = 198973;
16'd6450 : result1 = 197345;
16'd6656 : result1 = 289682;
16'd6657 : result1 = 285117;
16'd6658 : result1 = 281125;
16'd6659 : result1 = 277556;
16'd6660 : result1 = 274316;
16'd6661 : result1 = 271336;
16'd6662 : result1 = 268570;
16'd6663 : result1 = 265982;
16'd6664 : result1 = 263543;
16'd6665 : result1 = 261232;
16'd6666 : result1 = 259032;
16'd6667 : result1 = 256927;
16'd6668 : result1 = 254906;
16'd6669 : result1 = 252959;
16'd6670 : result1 = 251077;
16'd6671 : result1 = 249253;
16'd6672 : result1 = 247480;
16'd6673 : result1 = 245753;
16'd6674 : result1 = 244067;
16'd6675 : result1 = 242417;
16'd6676 : result1 = 240801;
16'd6677 : result1 = 239213;
16'd6678 : result1 = 237652;
16'd6679 : result1 = 236115;
16'd6680 : result1 = 234597;
16'd6681 : result1 = 233099;
16'd6682 : result1 = 231616;
16'd6683 : result1 = 230148;
16'd6684 : result1 = 228691;
16'd6685 : result1 = 227245;
16'd6686 : result1 = 225808;
16'd6687 : result1 = 224377;
16'd6688 : result1 = 222951;
16'd6689 : result1 = 221530;
16'd6690 : result1 = 220110;
16'd6691 : result1 = 218691;
16'd6692 : result1 = 217271;
16'd6693 : result1 = 215850;
16'd6694 : result1 = 214424;
16'd6695 : result1 = 212993;
16'd6696 : result1 = 211554;
16'd6697 : result1 = 210108;
16'd6698 : result1 = 208651;
16'd6699 : result1 = 207182;
16'd6700 : result1 = 205699;
16'd6701 : result1 = 204199;
16'd6702 : result1 = 202682;
16'd6703 : result1 = 201144;
16'd6704 : result1 = 199582;
16'd6705 : result1 = 197994;
16'd6706 : result1 = 196376;
16'd6912 : result1 = 285902;
16'd6913 : result1 = 281641;
16'd6914 : result1 = 277888;
16'd6915 : result1 = 274517;
16'd6916 : result1 = 271443;
16'd6917 : result1 = 268608;
16'd6918 : result1 = 265969;
16'd6919 : result1 = 263494;
16'd6920 : result1 = 261157;
16'd6921 : result1 = 258938;
16'd6922 : result1 = 256821;
16'd6923 : result1 = 254794;
16'd6924 : result1 = 252844;
16'd6925 : result1 = 250962;
16'd6926 : result1 = 249141;
16'd6927 : result1 = 247374;
16'd6928 : result1 = 245654;
16'd6929 : result1 = 243977;
16'd6930 : result1 = 242338;
16'd6931 : result1 = 240733;
16'd6932 : result1 = 239158;
16'd6933 : result1 = 237610;
16'd6934 : result1 = 236086;
16'd6935 : result1 = 234584;
16'd6936 : result1 = 233101;
16'd6937 : result1 = 231634;
16'd6938 : result1 = 230182;
16'd6939 : result1 = 228743;
16'd6940 : result1 = 227314;
16'd6941 : result1 = 225894;
16'd6942 : result1 = 224482;
16'd6943 : result1 = 223076;
16'd6944 : result1 = 221674;
16'd6945 : result1 = 220274;
16'd6946 : result1 = 218876;
16'd6947 : result1 = 217478;
16'd6948 : result1 = 216078;
16'd6949 : result1 = 214675;
16'd6950 : result1 = 213267;
16'd6951 : result1 = 211853;
16'd6952 : result1 = 210432;
16'd6953 : result1 = 209001;
16'd6954 : result1 = 207559;
16'd6955 : result1 = 206105;
16'd6956 : result1 = 204636;
16'd6957 : result1 = 203151;
16'd6958 : result1 = 201646;
16'd6959 : result1 = 200120;
16'd6960 : result1 = 198570;
16'd6961 : result1 = 196993;
16'd6962 : result1 = 195386;
16'd7168 : result1 = 282037;
16'd7169 : result1 = 278084;
16'd7170 : result1 = 274577;
16'd7171 : result1 = 271409;
16'd7172 : result1 = 268507;
16'd7173 : result1 = 265822;
16'd7174 : result1 = 263314;
16'd7175 : result1 = 260955;
16'd7176 : result1 = 258722;
16'd7177 : result1 = 256598;
16'd7178 : result1 = 254568;
16'd7179 : result1 = 252619;
16'd7180 : result1 = 250742;
16'd7181 : result1 = 248928;
16'd7182 : result1 = 247170;
16'd7183 : result1 = 245461;
16'd7184 : result1 = 243796;
16'd7185 : result1 = 242170;
16'd7186 : result1 = 240579;
16'd7187 : result1 = 239019;
16'd7188 : result1 = 237487;
16'd7189 : result1 = 235979;
16'd7190 : result1 = 234494;
16'd7191 : result1 = 233027;
16'd7192 : result1 = 231578;
16'd7193 : result1 = 230144;
16'd7194 : result1 = 228724;
16'd7195 : result1 = 227314;
16'd7196 : result1 = 225913;
16'd7197 : result1 = 224521;
16'd7198 : result1 = 223134;
16'd7199 : result1 = 221753;
16'd7200 : result1 = 220374;
16'd7201 : result1 = 218997;
16'd7202 : result1 = 217621;
16'd7203 : result1 = 216243;
16'd7204 : result1 = 214863;
16'd7205 : result1 = 213479;
16'd7206 : result1 = 212090;
16'd7207 : result1 = 210693;
16'd7208 : result1 = 209289;
16'd7209 : result1 = 207874;
16'd7210 : result1 = 206448;
16'd7211 : result1 = 205009;
16'd7212 : result1 = 203554;
16'd7213 : result1 = 202082;
16'd7214 : result1 = 200590;
16'd7215 : result1 = 199076;
16'd7216 : result1 = 197538;
16'd7217 : result1 = 195972;
16'd7218 : result1 = 194375;
16'd7424 : result1 = 278115;
16'd7425 : result1 = 274469;
16'd7426 : result1 = 271209;
16'd7427 : result1 = 268246;
16'd7428 : result1 = 265520;
16'd7429 : result1 = 262986;
16'd7430 : result1 = 260612;
16'd7431 : result1 = 258372;
16'd7432 : result1 = 256246;
16'd7433 : result1 = 254219;
16'd7434 : result1 = 252277;
16'd7435 : result1 = 250409;
16'd7436 : result1 = 248607;
16'd7437 : result1 = 246861;
16'd7438 : result1 = 245167;
16'd7439 : result1 = 243517;
16'd7440 : result1 = 241908;
16'd7441 : result1 = 240334;
16'd7442 : result1 = 238792;
16'd7443 : result1 = 237278;
16'd7444 : result1 = 235789;
16'd7445 : result1 = 234323;
16'd7446 : result1 = 232876;
16'd7447 : result1 = 231446;
16'd7448 : result1 = 230032;
16'd7449 : result1 = 228632;
16'd7450 : result1 = 227242;
16'd7451 : result1 = 225862;
16'd7452 : result1 = 224491;
16'd7453 : result1 = 223125;
16'd7454 : result1 = 221765;
16'd7455 : result1 = 220408;
16'd7456 : result1 = 219054;
16'd7457 : result1 = 217700;
16'd7458 : result1 = 216345;
16'd7459 : result1 = 214988;
16'd7460 : result1 = 213628;
16'd7461 : result1 = 212264;
16'd7462 : result1 = 210893;
16'd7463 : result1 = 209514;
16'd7464 : result1 = 208126;
16'd7465 : result1 = 206728;
16'd7466 : result1 = 205317;
16'd7467 : result1 = 203893;
16'd7468 : result1 = 202452;
16'd7469 : result1 = 200993;
16'd7470 : result1 = 199514;
16'd7471 : result1 = 198013;
16'd7472 : result1 = 196486;
16'd7473 : result1 = 194931;
16'd7474 : result1 = 193344;
16'd7680 : result1 = 274160;
16'd7681 : result1 = 270816;
16'd7682 : result1 = 267801;
16'd7683 : result1 = 265043;
16'd7684 : result1 = 262493;
16'd7685 : result1 = 260112;
16'd7686 : result1 = 257872;
16'd7687 : result1 = 255753;
16'd7688 : result1 = 253735;
16'd7689 : result1 = 251806;
16'd7690 : result1 = 249954;
16'd7691 : result1 = 248168;
16'd7692 : result1 = 246441;
16'd7693 : result1 = 244765;
16'd7694 : result1 = 243135;
16'd7695 : result1 = 241546;
16'd7696 : result1 = 239993;
16'd7697 : result1 = 238472;
16'd7698 : result1 = 236979;
16'd7699 : result1 = 235512;
16'd7700 : result1 = 234067;
16'd7701 : result1 = 232642;
16'd7702 : result1 = 231235;
16'd7703 : result1 = 229843;
16'd7704 : result1 = 228464;
16'd7705 : result1 = 227097;
16'd7706 : result1 = 225739;
16'd7707 : result1 = 224390;
16'd7708 : result1 = 223047;
16'd7709 : result1 = 221709;
16'd7710 : result1 = 220375;
16'd7711 : result1 = 219044;
16'd7712 : result1 = 217713;
16'd7713 : result1 = 216382;
16'd7714 : result1 = 215050;
16'd7715 : result1 = 213714;
16'd7716 : result1 = 212374;
16'd7717 : result1 = 211029;
16'd7718 : result1 = 209676;
16'd7719 : result1 = 208315;
16'd7720 : result1 = 206945;
16'd7721 : result1 = 205563;
16'd7722 : result1 = 204167;
16'd7723 : result1 = 202757;
16'd7724 : result1 = 201331;
16'd7725 : result1 = 199886;
16'd7726 : result1 = 198419;
16'd7727 : result1 = 196930;
16'd7728 : result1 = 195414;
16'd7729 : result1 = 193870;
16'd7730 : result1 = 192293;
16'd7936 : result1 = 270197;
16'd7937 : result1 = 267144;
16'd7938 : result1 = 264368;
16'd7939 : result1 = 261813;
16'd7940 : result1 = 259437;
16'd7941 : result1 = 257208;
16'd7942 : result1 = 255104;
16'd7943 : result1 = 253105;
16'd7944 : result1 = 251196;
16'd7945 : result1 = 249365;
16'd7946 : result1 = 247603;
16'd7947 : result1 = 245899;
16'd7948 : result1 = 244248;
16'd7949 : result1 = 242643;
16'd7950 : result1 = 241079;
16'd7951 : result1 = 239550;
16'd7952 : result1 = 238054;
16'd7953 : result1 = 236586;
16'd7954 : result1 = 235144;
16'd7955 : result1 = 233724;
16'd7956 : result1 = 232323;
16'd7957 : result1 = 230940;
16'd7958 : result1 = 229572;
16'd7959 : result1 = 228218;
16'd7960 : result1 = 226874;
16'd7961 : result1 = 225541;
16'd7962 : result1 = 224216;
16'd7963 : result1 = 222897;
16'd7964 : result1 = 221583;
16'd7965 : result1 = 220274;
16'd7966 : result1 = 218966;
16'd7967 : result1 = 217660;
16'd7968 : result1 = 216354;
16'd7969 : result1 = 215046;
16'd7970 : result1 = 213735;
16'd7971 : result1 = 212421;
16'd7972 : result1 = 211101;
16'd7973 : result1 = 209775;
16'd7974 : result1 = 208441;
16'd7975 : result1 = 207098;
16'd7976 : result1 = 205744;
16'd7977 : result1 = 204379;
16'd7978 : result1 = 202999;
16'd7979 : result1 = 201604;
16'd7980 : result1 = 200191;
16'd7981 : result1 = 198759;
16'd7982 : result1 = 197305;
16'd7983 : result1 = 195828;
16'd7984 : result1 = 194323;
16'd7985 : result1 = 192789;
16'd7986 : result1 = 191222;
16'd8192 : result1 = 266243;
16'd8193 : result1 = 263469;
16'd8194 : result1 = 260925;
16'd8195 : result1 = 258568;
16'd8196 : result1 = 256363;
16'd8197 : result1 = 254285;
16'd8198 : result1 = 252314;
16'd8199 : result1 = 250435;
16'd8200 : result1 = 248634;
16'd8201 : result1 = 246902;
16'd8202 : result1 = 245229;
16'd8203 : result1 = 243608;
16'd8204 : result1 = 242034;
16'd8205 : result1 = 240499;
16'd8206 : result1 = 239000;
16'd8207 : result1 = 237533;
16'd8208 : result1 = 236094;
16'd8209 : result1 = 234680;
16'd8210 : result1 = 233287;
16'd8211 : result1 = 231914;
16'd8212 : result1 = 230559;
16'd8213 : result1 = 229218;
16'd8214 : result1 = 227890;
16'd8215 : result1 = 226573;
16'd8216 : result1 = 225265;
16'd8217 : result1 = 223966;
16'd8218 : result1 = 222673;
16'd8219 : result1 = 221385;
16'd8220 : result1 = 220101;
16'd8221 : result1 = 218819;
16'd8222 : result1 = 217538;
16'd8223 : result1 = 216258;
16'd8224 : result1 = 214976;
16'd8225 : result1 = 213691;
16'd8226 : result1 = 212403;
16'd8227 : result1 = 211110;
16'd8228 : result1 = 209810;
16'd8229 : result1 = 208504;
16'd8230 : result1 = 207188;
16'd8231 : result1 = 205863;
16'd8232 : result1 = 204526;
16'd8233 : result1 = 203176;
16'd8234 : result1 = 201812;
16'd8235 : result1 = 200431;
16'd8236 : result1 = 199032;
16'd8237 : result1 = 197614;
16'd8238 : result1 = 196172;
16'd8239 : result1 = 194706;
16'd8240 : result1 = 193213;
16'd8241 : result1 = 191689;
16'd8242 : result1 = 190131;
16'd8448 : result1 = 262316;
16'd8449 : result1 = 259805;
16'd8450 : result1 = 257485;
16'd8451 : result1 = 255319;
16'd8452 : result1 = 253281;
16'd8453 : result1 = 251350;
16'd8454 : result1 = 249511;
16'd8455 : result1 = 247750;
16'd8456 : result1 = 246056;
16'd8457 : result1 = 244422;
16'd8458 : result1 = 242838;
16'd8459 : result1 = 241300;
16'd8460 : result1 = 239801;
16'd8461 : result1 = 238337;
16'd8462 : result1 = 236903;
16'd8463 : result1 = 235497;
16'd8464 : result1 = 234115;
16'd8465 : result1 = 232754;
16'd8466 : result1 = 231412;
16'd8467 : result1 = 230087;
16'd8468 : result1 = 228776;
16'd8469 : result1 = 227477;
16'd8470 : result1 = 226189;
16'd8471 : result1 = 224910;
16'd8472 : result1 = 223638;
16'd8473 : result1 = 222373;
16'd8474 : result1 = 221113;
16'd8475 : result1 = 219856;
16'd8476 : result1 = 218601;
16'd8477 : result1 = 217347;
16'd8478 : result1 = 216093;
16'd8479 : result1 = 214838;
16'd8480 : result1 = 213580;
16'd8481 : result1 = 212319;
16'd8482 : result1 = 211053;
16'd8483 : result1 = 209781;
16'd8484 : result1 = 208502;
16'd8485 : result1 = 207215;
16'd8486 : result1 = 205918;
16'd8487 : result1 = 204610;
16'd8488 : result1 = 203290;
16'd8489 : result1 = 201956;
16'd8490 : result1 = 200607;
16'd8491 : result1 = 199241;
16'd8492 : result1 = 197856;
16'd8493 : result1 = 196450;
16'd8494 : result1 = 195021;
16'd8495 : result1 = 193566;
16'd8496 : result1 = 192084;
16'd8497 : result1 = 190569;
16'd8498 : result1 = 189020;
16'd8704 : result1 = 258429;
16'd8705 : result1 = 256167;
16'd8706 : result1 = 254058;
16'd8707 : result1 = 252076;
16'd8708 : result1 = 250199;
16'd8709 : result1 = 248412;
16'd8710 : result1 = 246701;
16'd8711 : result1 = 245056;
16'd8712 : result1 = 243468;
16'd8713 : result1 = 241930;
16'd8714 : result1 = 240434;
16'd8715 : result1 = 238977;
16'd8716 : result1 = 237553;
16'd8717 : result1 = 236159;
16'd8718 : result1 = 234791;
16'd8719 : result1 = 233445;
16'd8720 : result1 = 232120;
16'd8721 : result1 = 230813;
16'd8722 : result1 = 229521;
16'd8723 : result1 = 228243;
16'd8724 : result1 = 226976;
16'd8725 : result1 = 225720;
16'd8726 : result1 = 224471;
16'd8727 : result1 = 223230;
16'd8728 : result1 = 221995;
16'd8729 : result1 = 220764;
16'd8730 : result1 = 219536;
16'd8731 : result1 = 218309;
16'd8732 : result1 = 217084;
16'd8733 : result1 = 215858;
16'd8734 : result1 = 214631;
16'd8735 : result1 = 213401;
16'd8736 : result1 = 212168;
16'd8737 : result1 = 210930;
16'd8738 : result1 = 209686;
16'd8739 : result1 = 208435;
16'd8740 : result1 = 207177;
16'd8741 : result1 = 205909;
16'd8742 : result1 = 204630;
16'd8743 : result1 = 203340;
16'd8744 : result1 = 202037;
16'd8745 : result1 = 200719;
16'd8746 : result1 = 199385;
16'd8747 : result1 = 198033;
16'd8748 : result1 = 196662;
16'd8749 : result1 = 195269;
16'd8750 : result1 = 193852;
16'd8751 : result1 = 192408;
16'd8752 : result1 = 190935;
16'd8753 : result1 = 189430;
16'd8754 : result1 = 187890;
16'd8960 : result1 = 254594;
16'd8961 : result1 = 252564;
16'd8962 : result1 = 250655;
16'd8963 : result1 = 248848;
16'd8964 : result1 = 247127;
16'd8965 : result1 = 245478;
16'd8966 : result1 = 243892;
16'd8967 : result1 = 242360;
16'd8968 : result1 = 240875;
16'd8969 : result1 = 239430;
16'd8970 : result1 = 238022;
16'd8971 : result1 = 236645;
16'd8972 : result1 = 235295;
16'd8973 : result1 = 233970;
16'd8974 : result1 = 232666;
16'd8975 : result1 = 231381;
16'd8976 : result1 = 230112;
16'd8977 : result1 = 228858;
16'd8978 : result1 = 227616;
16'd8979 : result1 = 226384;
16'd8980 : result1 = 225162;
16'd8981 : result1 = 223948;
16'd8982 : result1 = 222739;
16'd8983 : result1 = 221536;
16'd8984 : result1 = 220336;
16'd8985 : result1 = 219139;
16'd8986 : result1 = 217943;
16'd8987 : result1 = 216748;
16'd8988 : result1 = 215552;
16'd8989 : result1 = 214354;
16'd8990 : result1 = 213153;
16'd8991 : result1 = 211949;
16'd8992 : result1 = 210740;
16'd8993 : result1 = 209525;
16'd8994 : result1 = 208303;
16'd8995 : result1 = 207074;
16'd8996 : result1 = 205835;
16'd8997 : result1 = 204587;
16'd8998 : result1 = 203327;
16'd8999 : result1 = 202054;
16'd9000 : result1 = 200767;
16'd9001 : result1 = 199465;
16'd9002 : result1 = 198146;
16'd9003 : result1 = 196808;
16'd9004 : result1 = 195450;
16'd9005 : result1 = 194070;
16'd9006 : result1 = 192664;
16'd9007 : result1 = 191231;
16'd9008 : result1 = 189769;
16'd9009 : result1 = 188273;
16'd9010 : result1 = 186740;
16'd9216 : result1 = 250820;
16'd9217 : result1 = 249005;
16'd9218 : result1 = 247284;
16'd9219 : result1 = 245644;
16'd9220 : result1 = 244070;
16'd9221 : result1 = 242555;
16'd9222 : result1 = 241089;
16'd9223 : result1 = 239666;
16'd9224 : result1 = 238281;
16'd9225 : result1 = 236929;
16'd9226 : result1 = 235605;
16'd9227 : result1 = 234306;
16'd9228 : result1 = 233030;
16'd9229 : result1 = 231772;
16'd9230 : result1 = 230532;
16'd9231 : result1 = 229306;
16'd9232 : result1 = 228093;
16'd9233 : result1 = 226891;
16'd9234 : result1 = 225698;
16'd9235 : result1 = 224514;
16'd9236 : result1 = 223336;
16'd9237 : result1 = 222163;
16'd9238 : result1 = 220994;
16'd9239 : result1 = 219828;
16'd9240 : result1 = 218663;
16'd9241 : result1 = 217500;
16'd9242 : result1 = 216336;
16'd9243 : result1 = 215172;
16'd9244 : result1 = 214005;
16'd9245 : result1 = 212835;
16'd9246 : result1 = 211661;
16'd9247 : result1 = 210482;
16'd9248 : result1 = 209297;
16'd9249 : result1 = 208105;
16'd9250 : result1 = 206905;
16'd9251 : result1 = 205697;
16'd9252 : result1 = 204478;
16'd9253 : result1 = 203249;
16'd9254 : result1 = 202007;
16'd9255 : result1 = 200751;
16'd9256 : result1 = 199481;
16'd9257 : result1 = 198195;
16'd9258 : result1 = 196890;
16'd9259 : result1 = 195567;
16'd9260 : result1 = 194222;
16'd9261 : result1 = 192853;
16'd9262 : result1 = 191459;
16'd9263 : result1 = 190037;
16'd9264 : result1 = 188584;
16'd9265 : result1 = 187096;
16'd9266 : result1 = 185571;
16'd9472 : result1 = 247112;
16'd9473 : result1 = 245497;
16'd9474 : result1 = 243953;
16'd9475 : result1 = 242469;
16'd9476 : result1 = 241036;
16'd9477 : result1 = 239647;
16'd9478 : result1 = 238297;
16'd9479 : result1 = 236980;
16'd9480 : result1 = 235692;
16'd9481 : result1 = 234428;
16'd9482 : result1 = 233187;
16'd9483 : result1 = 231965;
16'd9484 : result1 = 230760;
16'd9485 : result1 = 229569;
16'd9486 : result1 = 228391;
16'd9487 : result1 = 227224;
16'd9488 : result1 = 226066;
16'd9489 : result1 = 224915;
16'd9490 : result1 = 223771;
16'd9491 : result1 = 222633;
16'd9492 : result1 = 221498;
16'd9493 : result1 = 220366;
16'd9494 : result1 = 219236;
16'd9495 : result1 = 218107;
16'd9496 : result1 = 216978;
16'd9497 : result1 = 215848;
16'd9498 : result1 = 214717;
16'd9499 : result1 = 213582;
16'd9500 : result1 = 212444;
16'd9501 : result1 = 211302;
16'd9502 : result1 = 210154;
16'd9503 : result1 = 209001;
16'd9504 : result1 = 207840;
16'd9505 : result1 = 206671;
16'd9506 : result1 = 205493;
16'd9507 : result1 = 204305;
16'd9508 : result1 = 203106;
16'd9509 : result1 = 201896;
16'd9510 : result1 = 200672;
16'd9511 : result1 = 199433;
16'd9512 : result1 = 198179;
16'd9513 : result1 = 196908;
16'd9514 : result1 = 195619;
16'd9515 : result1 = 194308;
16'd9516 : result1 = 192976;
16'd9517 : result1 = 191620;
16'd9518 : result1 = 190237;
16'd9519 : result1 = 188825;
16'd9520 : result1 = 187381;
16'd9521 : result1 = 185901;
16'd9522 : result1 = 184383;
16'd9728 : result1 = 243478;
16'd9729 : result1 = 242047;
16'd9730 : result1 = 240666;
16'd9731 : result1 = 239329;
16'd9732 : result1 = 238029;
16'd9733 : result1 = 236762;
16'd9734 : result1 = 235522;
16'd9735 : result1 = 234306;
16'd9736 : result1 = 233111;
16'd9737 : result1 = 231934;
16'd9738 : result1 = 230773;
16'd9739 : result1 = 229625;
16'd9740 : result1 = 228489;
16'd9741 : result1 = 227363;
16'd9742 : result1 = 226246;
16'd9743 : result1 = 225136;
16'd9744 : result1 = 224032;
16'd9745 : result1 = 222932;
16'd9746 : result1 = 221836;
16'd9747 : result1 = 220743;
16'd9748 : result1 = 219651;
16'd9749 : result1 = 218560;
16'd9750 : result1 = 217468;
16'd9751 : result1 = 216376;
16'd9752 : result1 = 215282;
16'd9753 : result1 = 214185;
16'd9754 : result1 = 213085;
16'd9755 : result1 = 211981;
16'd9756 : result1 = 210872;
16'd9757 : result1 = 209757;
16'd9758 : result1 = 208635;
16'd9759 : result1 = 207506;
16'd9760 : result1 = 206369;
16'd9761 : result1 = 205223;
16'd9762 : result1 = 204066;
16'd9763 : result1 = 202899;
16'd9764 : result1 = 201720;
16'd9765 : result1 = 200528;
16'd9766 : result1 = 199322;
16'd9767 : result1 = 198100;
16'd9768 : result1 = 196862;
16'd9769 : result1 = 195606;
16'd9770 : result1 = 194331;
16'd9771 : result1 = 193034;
16'd9772 : result1 = 191714;
16'd9773 : result1 = 190369;
16'd9774 : result1 = 188997;
16'd9775 : result1 = 187595;
16'd9776 : result1 = 186159;
16'd9777 : result1 = 184688;
16'd9778 : result1 = 183176;
16'd9984 : result1 = 239919;
16'd9985 : result1 = 238657;
16'd9986 : result1 = 237429;
16'd9987 : result1 = 236229;
16'd9988 : result1 = 235055;
16'd9989 : result1 = 233901;
16'd9990 : result1 = 232766;
16'd9991 : result1 = 231647;
16'd9992 : result1 = 230542;
16'd9993 : result1 = 229448;
16'd9994 : result1 = 228364;
16'd9995 : result1 = 227288;
16'd9996 : result1 = 226220;
16'd9997 : result1 = 225158;
16'd9998 : result1 = 224100;
16'd9999 : result1 = 223045;
16'd10000 : result1 = 221994;
16'd10001 : result1 = 220944;
16'd10002 : result1 = 219895;
16'd10003 : result1 = 218846;
16'd10004 : result1 = 217796;
16'd10005 : result1 = 216745;
16'd10006 : result1 = 215692;
16'd10007 : result1 = 214636;
16'd10008 : result1 = 213576;
16'd10009 : result1 = 212512;
16'd10010 : result1 = 211443;
16'd10011 : result1 = 210368;
16'd10012 : result1 = 209287;
16'd10013 : result1 = 208199;
16'd10014 : result1 = 207103;
16'd10015 : result1 = 205999;
16'd10016 : result1 = 204885;
16'd10017 : result1 = 203761;
16'd10018 : result1 = 202626;
16'd10019 : result1 = 201480;
16'd10020 : result1 = 200320;
16'd10021 : result1 = 199146;
16'd10022 : result1 = 197958;
16'd10023 : result1 = 196753;
16'd10024 : result1 = 195530;
16'd10025 : result1 = 194289;
16'd10026 : result1 = 193028;
16'd10027 : result1 = 191744;
16'd10028 : result1 = 190436;
16'd10029 : result1 = 189102;
16'd10030 : result1 = 187740;
16'd10031 : result1 = 186347;
16'd10032 : result1 = 184920;
16'd10033 : result1 = 183456;
16'd10034 : result1 = 181950;
16'd10240 : result1 = 236439;
16'd10241 : result1 = 235332;
16'd10242 : result1 = 234244;
16'd10243 : result1 = 233173;
16'd10244 : result1 = 232116;
16'd10245 : result1 = 231070;
16'd10246 : result1 = 230035;
16'd10247 : result1 = 229008;
16'd10248 : result1 = 227988;
16'd10249 : result1 = 226974;
16'd10250 : result1 = 225964;
16'd10251 : result1 = 224958;
16'd10252 : result1 = 223955;
16'd10253 : result1 = 222954;
16'd10254 : result1 = 221954;
16'd10255 : result1 = 220954;
16'd10256 : result1 = 219953;
16'd10257 : result1 = 218952;
16'd10258 : result1 = 217949;
16'd10259 : result1 = 216944;
16'd10260 : result1 = 215935;
16'd10261 : result1 = 214923;
16'd10262 : result1 = 213908;
16'd10263 : result1 = 212887;
16'd10264 : result1 = 211861;
16'd10265 : result1 = 210829;
16'd10266 : result1 = 209791;
16'd10267 : result1 = 208745;
16'd10268 : result1 = 207692;
16'd10269 : result1 = 206631;
16'd10270 : result1 = 205561;
16'd10271 : result1 = 204480;
16'd10272 : result1 = 203390;
16'd10273 : result1 = 202288;
16'd10274 : result1 = 201174;
16'd10275 : result1 = 200047;
16'd10276 : result1 = 198906;
16'd10277 : result1 = 197751;
16'd10278 : result1 = 196579;
16'd10279 : result1 = 195391;
16'd10280 : result1 = 194184;
16'd10281 : result1 = 192957;
16'd10282 : result1 = 191709;
16'd10283 : result1 = 190438;
16'd10284 : result1 = 189142;
16'd10285 : result1 = 187819;
16'd10286 : result1 = 186467;
16'd10287 : result1 = 185083;
16'd10288 : result1 = 183663;
16'd10289 : result1 = 182205;
16'd10290 : result1 = 180704;
16'd10496 : result1 = 233039;
16'd10497 : result1 = 232074;
16'd10498 : result1 = 231116;
16'd10499 : result1 = 230163;
16'd10500 : result1 = 229216;
16'd10501 : result1 = 228271;
16'd10502 : result1 = 227330;
16'd10503 : result1 = 226390;
16'd10504 : result1 = 225452;
16'd10505 : result1 = 224514;
16'd10506 : result1 = 223576;
16'd10507 : result1 = 222637;
16'd10508 : result1 = 221697;
16'd10509 : result1 = 220755;
16'd10510 : result1 = 219810;
16'd10511 : result1 = 218863;
16'd10512 : result1 = 217913;
16'd10513 : result1 = 216959;
16'd10514 : result1 = 216001;
16'd10515 : result1 = 215038;
16'd10516 : result1 = 214070;
16'd10517 : result1 = 213096;
16'd10518 : result1 = 212117;
16'd10519 : result1 = 211131;
16'd10520 : result1 = 210138;
16'd10521 : result1 = 209138;
16'd10522 : result1 = 208130;
16'd10523 : result1 = 207113;
16'd10524 : result1 = 206088;
16'd10525 : result1 = 205052;
16'd10526 : result1 = 204007;
16'd10527 : result1 = 202951;
16'd10528 : result1 = 201883;
16'd10529 : result1 = 200803;
16'd10530 : result1 = 199709;
16'd10531 : result1 = 198602;
16'd10532 : result1 = 197480;
16'd10533 : result1 = 196342;
16'd10534 : result1 = 195188;
16'd10535 : result1 = 194015;
16'd10536 : result1 = 192823;
16'd10537 : result1 = 191611;
16'd10538 : result1 = 190376;
16'd10539 : result1 = 189117;
16'd10540 : result1 = 187832;
16'd10541 : result1 = 186520;
16'd10542 : result1 = 185177;
16'd10543 : result1 = 183801;
16'd10544 : result1 = 182388;
16'd10545 : result1 = 180936;
16'd10546 : result1 = 179440;
16'd10752 : result1 = 229719;
16'd10753 : result1 = 228883;
16'd10754 : result1 = 228044;
16'd10755 : result1 = 227202;
16'd10756 : result1 = 226357;
16'd10757 : result1 = 225508;
16'd10758 : result1 = 224655;
16'd10759 : result1 = 223798;
16'd10760 : result1 = 222937;
16'd10761 : result1 = 222071;
16'd10762 : result1 = 221201;
16'd10763 : result1 = 220326;
16'd10764 : result1 = 219447;
16'd10765 : result1 = 218562;
16'd10766 : result1 = 217671;
16'd10767 : result1 = 216775;
16'd10768 : result1 = 215873;
16'd10769 : result1 = 214965;
16'd10770 : result1 = 214051;
16'd10771 : result1 = 213129;
16'd10772 : result1 = 212201;
16'd10773 : result1 = 211265;
16'd10774 : result1 = 210321;
16'd10775 : result1 = 209369;
16'd10776 : result1 = 208409;
16'd10777 : result1 = 207440;
16'd10778 : result1 = 206461;
16'd10779 : result1 = 205473;
16'd10780 : result1 = 204474;
16'd10781 : result1 = 203465;
16'd10782 : result1 = 202444;
16'd10783 : result1 = 201411;
16'd10784 : result1 = 200365;
16'd10785 : result1 = 199306;
16'd10786 : result1 = 198233;
16'd10787 : result1 = 197145;
16'd10788 : result1 = 196042;
16'd10789 : result1 = 194921;
16'd10790 : result1 = 193783;
16'd10791 : result1 = 192626;
16'd10792 : result1 = 191449;
16'd10793 : result1 = 190250;
16'd10794 : result1 = 189028;
16'd10795 : result1 = 187781;
16'd10796 : result1 = 186507;
16'd10797 : result1 = 185204;
16'd10798 : result1 = 183870;
16'd10799 : result1 = 182501;
16'd10800 : result1 = 181095;
16'd10801 : result1 = 179648;
16'd10802 : result1 = 178156;
16'd11008 : result1 = 226478;
16'd11009 : result1 = 225760;
16'd11010 : result1 = 225031;
16'd11011 : result1 = 224291;
16'd11012 : result1 = 223541;
16'd11013 : result1 = 222780;
16'd11014 : result1 = 222010;
16'd11015 : result1 = 221231;
16'd11016 : result1 = 220444;
16'd11017 : result1 = 219647;
16'd11018 : result1 = 218842;
16'd11019 : result1 = 218029;
16'd11020 : result1 = 217207;
16'd11021 : result1 = 216377;
16'd11022 : result1 = 215539;
16'd11023 : result1 = 214692;
16'd11024 : result1 = 213837;
16'd11025 : result1 = 212973;
16'd11026 : result1 = 212101;
16'd11027 : result1 = 211220;
16'd11028 : result1 = 210330;
16'd11029 : result1 = 209430;
16'd11030 : result1 = 208521;
16'd11031 : result1 = 207603;
16'd11032 : result1 = 206674;
16'd11033 : result1 = 205735;
16'd11034 : result1 = 204785;
16'd11035 : result1 = 203825;
16'd11036 : result1 = 202852;
16'd11037 : result1 = 201868;
16'd11038 : result1 = 200871;
16'd11039 : result1 = 199861;
16'd11040 : result1 = 198837;
16'd11041 : result1 = 197799;
16'd11042 : result1 = 196746;
16'd11043 : result1 = 195677;
16'd11044 : result1 = 194591;
16'd11045 : result1 = 193488;
16'd11046 : result1 = 192366;
16'd11047 : result1 = 191224;
16'd11048 : result1 = 190061;
16'd11049 : result1 = 188875;
16'd11050 : result1 = 187665;
16'd11051 : result1 = 186429;
16'd11052 : result1 = 185166;
16'd11053 : result1 = 183872;
16'd11054 : result1 = 182546;
16'd11055 : result1 = 181185;
16'd11056 : result1 = 179785;
16'd11057 : result1 = 178342;
16'd11058 : result1 = 176852;
16'd11264 : result1 = 223316;
16'd11265 : result1 = 222706;
16'd11266 : result1 = 222077;
16'd11267 : result1 = 221431;
16'd11268 : result1 = 220769;
16'd11269 : result1 = 220091;
16'd11270 : result1 = 219399;
16'd11271 : result1 = 218694;
16'd11272 : result1 = 217975;
16'd11273 : result1 = 217244;
16'd11274 : result1 = 216501;
16'd11275 : result1 = 215746;
16'd11276 : result1 = 214980;
16'd11277 : result1 = 214202;
16'd11278 : result1 = 213414;
16'd11279 : result1 = 212615;
16'd11280 : result1 = 211805;
16'd11281 : result1 = 210984;
16'd11282 : result1 = 210152;
16'd11283 : result1 = 209310;
16'd11284 : result1 = 208457;
16'd11285 : result1 = 207593;
16'd11286 : result1 = 206718;
16'd11287 : result1 = 205832;
16'd11288 : result1 = 204935;
16'd11289 : result1 = 204025;
16'd11290 : result1 = 203104;
16'd11291 : result1 = 202170;
16'd11292 : result1 = 201223;
16'd11293 : result1 = 200263;
16'd11294 : result1 = 199290;
16'd11295 : result1 = 198302;
16'd11296 : result1 = 197300;
16'd11297 : result1 = 196282;
16'd11298 : result1 = 195248;
16'd11299 : result1 = 194198;
16'd11300 : result1 = 193130;
16'd11301 : result1 = 192043;
16'd11302 : result1 = 190936;
16'd11303 : result1 = 189809;
16'd11304 : result1 = 188659;
16'd11305 : result1 = 187486;
16'd11306 : result1 = 186288;
16'd11307 : result1 = 185063;
16'd11308 : result1 = 183810;
16'd11309 : result1 = 182525;
16'd11310 : result1 = 181206;
16'd11311 : result1 = 179851;
16'd11312 : result1 = 178456;
16'd11313 : result1 = 177017;
16'd11314 : result1 = 175529;
16'd11520 : result1 = 220232;
16'd11521 : result1 = 219719;
16'd11522 : result1 = 219182;
16'd11523 : result1 = 218622;
16'd11524 : result1 = 218042;
16'd11525 : result1 = 217441;
16'd11526 : result1 = 216822;
16'd11527 : result1 = 216185;
16'd11528 : result1 = 215532;
16'd11529 : result1 = 214862;
16'd11530 : result1 = 214178;
16'd11531 : result1 = 213479;
16'd11532 : result1 = 212765;
16'd11533 : result1 = 212038;
16'd11534 : result1 = 211298;
16'd11535 : result1 = 210544;
16'd11536 : result1 = 209778;
16'd11537 : result1 = 208998;
16'd11538 : result1 = 208206;
16'd11539 : result1 = 207402;
16'd11540 : result1 = 206585;
16'd11541 : result1 = 205756;
16'd11542 : result1 = 204914;
16'd11543 : result1 = 204059;
16'd11544 : result1 = 203191;
16'd11545 : result1 = 202310;
16'd11546 : result1 = 201416;
16'd11547 : result1 = 200509;
16'd11548 : result1 = 199587;
16'd11549 : result1 = 198651;
16'd11550 : result1 = 197701;
16'd11551 : result1 = 196735;
16'd11552 : result1 = 195753;
16'd11553 : result1 = 194756;
16'd11554 : result1 = 193741;
16'd11555 : result1 = 192708;
16'd11556 : result1 = 191657;
16'd11557 : result1 = 190586;
16'd11558 : result1 = 189494;
16'd11559 : result1 = 188381;
16'd11560 : result1 = 187245;
16'd11561 : result1 = 186084;
16'd11562 : result1 = 184897;
16'd11563 : result1 = 183683;
16'd11564 : result1 = 182438;
16'd11565 : result1 = 181161;
16'd11566 : result1 = 179850;
16'd11567 : result1 = 178500;
16'd11568 : result1 = 177109;
16'd11569 : result1 = 175673;
16'd11570 : result1 = 174185;
16'd11776 : result1 = 217223;
16'd11777 : result1 = 216799;
16'd11778 : result1 = 216346;
16'd11779 : result1 = 215865;
16'd11780 : result1 = 215360;
16'd11781 : result1 = 214831;
16'd11782 : result1 = 214279;
16'd11783 : result1 = 213707;
16'd11784 : result1 = 213115;
16'd11785 : result1 = 212504;
16'd11786 : result1 = 211875;
16'd11787 : result1 = 211229;
16'd11788 : result1 = 210566;
16'd11789 : result1 = 209887;
16'd11790 : result1 = 209192;
16'd11791 : result1 = 208482;
16'd11792 : result1 = 207757;
16'd11793 : result1 = 207018;
16'd11794 : result1 = 206264;
16'd11795 : result1 = 205496;
16'd11796 : result1 = 204714;
16'd11797 : result1 = 203918;
16'd11798 : result1 = 203107;
16'd11799 : result1 = 202283;
16'd11800 : result1 = 201445;
16'd11801 : result1 = 200592;
16'd11802 : result1 = 199724;
16'd11803 : result1 = 198842;
16'd11804 : result1 = 197945;
16'd11805 : result1 = 197033;
16'd11806 : result1 = 196104;
16'd11807 : result1 = 195160;
16'd11808 : result1 = 194198;
16'd11809 : result1 = 193220;
16'd11810 : result1 = 192223;
16'd11811 : result1 = 191208;
16'd11812 : result1 = 190173;
16'd11813 : result1 = 189117;
16'd11814 : result1 = 188041;
16'd11815 : result1 = 186941;
16'd11816 : result1 = 185817;
16'd11817 : result1 = 184668;
16'd11818 : result1 = 183492;
16'd11819 : result1 = 182287;
16'd11820 : result1 = 181051;
16'd11821 : result1 = 179782;
16'd11822 : result1 = 178477;
16'd11823 : result1 = 177132;
16'd11824 : result1 = 175744;
16'd11825 : result1 = 174309;
16'd11826 : result1 = 172822;
16'd12032 : result1 = 214288;
16'd12033 : result1 = 213944;
16'd12034 : result1 = 213567;
16'd12035 : result1 = 213159;
16'd12036 : result1 = 212723;
16'd12037 : result1 = 212261;
16'd12038 : result1 = 211773;
16'd12039 : result1 = 211261;
16'd12040 : result1 = 210726;
16'd12041 : result1 = 210170;
16'd12042 : result1 = 209593;
16'd12043 : result1 = 208997;
16'd12044 : result1 = 208382;
16'd12045 : result1 = 207748;
16'd12046 : result1 = 207097;
16'd12047 : result1 = 206429;
16'd12048 : result1 = 205744;
16'd12049 : result1 = 205043;
16'd12050 : result1 = 204326;
16'd12051 : result1 = 203593;
16'd12052 : result1 = 202844;
16'd12053 : result1 = 202080;
16'd12054 : result1 = 201301;
16'd12055 : result1 = 200506;
16'd12056 : result1 = 199696;
16'd12057 : result1 = 198870;
16'd12058 : result1 = 198028;
16'd12059 : result1 = 197171;
16'd12060 : result1 = 196298;
16'd12061 : result1 = 195408;
16'd12062 : result1 = 194501;
16'd12063 : result1 = 193577;
16'd12064 : result1 = 192635;
16'd12065 : result1 = 191675;
16'd12066 : result1 = 190696;
16'd12067 : result1 = 189698;
16'd12068 : result1 = 188679;
16'd12069 : result1 = 187638;
16'd12070 : result1 = 186575;
16'd12071 : result1 = 185489;
16'd12072 : result1 = 184377;
16'd12073 : result1 = 183239;
16'd12074 : result1 = 182073;
16'd12075 : result1 = 180878;
16'd12076 : result1 = 179649;
16'd12077 : result1 = 178387;
16'd12078 : result1 = 177087;
16'd12079 : result1 = 175746;
16'd12080 : result1 = 174360;
16'd12081 : result1 = 172926;
16'd12082 : result1 = 171437;
16'd12288 : result1 = 211424;
16'd12289 : result1 = 211152;
16'd12290 : result1 = 210845;
16'd12291 : result1 = 210504;
16'd12292 : result1 = 210132;
16'd12293 : result1 = 209731;
16'd12294 : result1 = 209301;
16'd12295 : result1 = 208845;
16'd12296 : result1 = 208365;
16'd12297 : result1 = 207860;
16'd12298 : result1 = 207333;
16'd12299 : result1 = 206784;
16'd12300 : result1 = 206214;
16'd12301 : result1 = 205624;
16'd12302 : result1 = 205014;
16'd12303 : result1 = 204386;
16'd12304 : result1 = 203739;
16'd12305 : result1 = 203075;
16'd12306 : result1 = 202393;
16'd12307 : result1 = 201694;
16'd12308 : result1 = 200977;
16'd12309 : result1 = 200244;
16'd12310 : result1 = 199495;
16'd12311 : result1 = 198728;
16'd12312 : result1 = 197945;
16'd12313 : result1 = 197145;
16'd12314 : result1 = 196329;
16'd12315 : result1 = 195496;
16'd12316 : result1 = 194645;
16'd12317 : result1 = 193777;
16'd12318 : result1 = 192891;
16'd12319 : result1 = 191987;
16'd12320 : result1 = 191064;
16'd12321 : result1 = 190122;
16'd12322 : result1 = 189161;
16'd12323 : result1 = 188178;
16'd12324 : result1 = 187174;
16'd12325 : result1 = 186148;
16'd12326 : result1 = 185099;
16'd12327 : result1 = 184025;
16'd12328 : result1 = 182925;
16'd12329 : result1 = 181797;
16'd12330 : result1 = 180641;
16'd12331 : result1 = 179453;
16'd12332 : result1 = 178232;
16'd12333 : result1 = 176975;
16'd12334 : result1 = 175680;
16'd12335 : result1 = 174342;
16'd12336 : result1 = 172958;
16'd12337 : result1 = 171523;
16'd12338 : result1 = 170031;
16'd12544 : result1 = 208628;
16'd12545 : result1 = 208422;
16'd12546 : result1 = 208179;
16'd12547 : result1 = 207899;
16'd12548 : result1 = 207586;
16'd12549 : result1 = 207241;
16'd12550 : result1 = 206866;
16'd12551 : result1 = 206462;
16'd12552 : result1 = 206032;
16'd12553 : result1 = 205575;
16'd12554 : result1 = 205095;
16'd12555 : result1 = 204590;
16'd12556 : result1 = 204063;
16'd12557 : result1 = 203514;
16'd12558 : result1 = 202944;
16'd12559 : result1 = 202354;
16'd12560 : result1 = 201744;
16'd12561 : result1 = 201114;
16'd12562 : result1 = 200466;
16'd12563 : result1 = 199799;
16'd12564 : result1 = 199114;
16'd12565 : result1 = 198410;
16'd12566 : result1 = 197689;
16'd12567 : result1 = 196950;
16'd12568 : result1 = 196193;
16'd12569 : result1 = 195419;
16'd12570 : result1 = 194626;
16'd12571 : result1 = 193816;
16'd12572 : result1 = 192988;
16'd12573 : result1 = 192141;
16'd12574 : result1 = 191275;
16'd12575 : result1 = 190390;
16'd12576 : result1 = 189486;
16'd12577 : result1 = 188561;
16'd12578 : result1 = 187616;
16'd12579 : result1 = 186649;
16'd12580 : result1 = 185660;
16'd12581 : result1 = 184648;
16'd12582 : result1 = 183611;
16'd12583 : result1 = 182549;
16'd12584 : result1 = 181459;
16'd12585 : result1 = 180342;
16'd12586 : result1 = 179194;
16'd12587 : result1 = 178014;
16'd12588 : result1 = 176799;
16'd12589 : result1 = 175547;
16'd12590 : result1 = 174255;
16'd12591 : result1 = 172919;
16'd12592 : result1 = 171536;
16'd12593 : result1 = 170099;
16'd12594 : result1 = 168603;
16'd12800 : result1 = 205899;
16'd12801 : result1 = 205753;
16'd12802 : result1 = 205566;
16'd12803 : result1 = 205342;
16'd12804 : result1 = 205083;
16'd12805 : result1 = 204790;
16'd12806 : result1 = 204466;
16'd12807 : result1 = 204111;
16'd12808 : result1 = 203727;
16'd12809 : result1 = 203316;
16'd12810 : result1 = 202879;
16'd12811 : result1 = 202416;
16'd12812 : result1 = 201930;
16'd12813 : result1 = 201420;
16'd12814 : result1 = 200887;
16'd12815 : result1 = 200333;
16'd12816 : result1 = 199758;
16'd12817 : result1 = 199161;
16'd12818 : result1 = 198545;
16'd12819 : result1 = 197909;
16'd12820 : result1 = 197253;
16'd12821 : result1 = 196579;
16'd12822 : result1 = 195885;
16'd12823 : result1 = 195172;
16'd12824 : result1 = 194441;
16'd12825 : result1 = 193691;
16'd12826 : result1 = 192921;
16'd12827 : result1 = 192133;
16'd12828 : result1 = 191326;
16'd12829 : result1 = 190500;
16'd12830 : result1 = 189654;
16'd12831 : result1 = 188787;
16'd12832 : result1 = 187901;
16'd12833 : result1 = 186993;
16'd12834 : result1 = 186063;
16'd12835 : result1 = 185111;
16'd12836 : result1 = 184136;
16'd12837 : result1 = 183137;
16'd12838 : result1 = 182112;
16'd12839 : result1 = 181061;
16'd12840 : result1 = 179982;
16'd12841 : result1 = 178873;
16'd12842 : result1 = 177733;
16'd12843 : result1 = 176560;
16'd12844 : result1 = 175351;
16'd12845 : result1 = 174103;
16'd12846 : result1 = 172813;
16'd12847 : result1 = 171478;
16'd12848 : result1 = 170094;
16'd12849 : result1 = 168653;
16'd12850 : result1 = 167152;
16'd13056 : result1 = 203233;
16'd13057 : result1 = 203140;
16'd13058 : result1 = 203006;
16'd13059 : result1 = 202833;
16'd13060 : result1 = 202624;
16'd13061 : result1 = 202379;
16'd13062 : result1 = 202101;
16'd13063 : result1 = 201791;
16'd13064 : result1 = 201451;
16'd13065 : result1 = 201082;
16'd13066 : result1 = 200686;
16'd13067 : result1 = 200263;
16'd13068 : result1 = 199814;
16'd13069 : result1 = 199341;
16'd13070 : result1 = 198844;
16'd13071 : result1 = 198324;
16'd13072 : result1 = 197781;
16'd13073 : result1 = 197217;
16'd13074 : result1 = 196631;
16'd13075 : result1 = 196025;
16'd13076 : result1 = 195398;
16'd13077 : result1 = 194750;
16'd13078 : result1 = 194083;
16'd13079 : result1 = 193395;
16'd13080 : result1 = 192688;
16'd13081 : result1 = 191961;
16'd13082 : result1 = 191214;
16'd13083 : result1 = 190448;
16'd13084 : result1 = 189661;
16'd13085 : result1 = 188854;
16'd13086 : result1 = 188027;
16'd13087 : result1 = 187178;
16'd13088 : result1 = 186308;
16'd13089 : result1 = 185416;
16'd13090 : result1 = 184502;
16'd13091 : result1 = 183564;
16'd13092 : result1 = 182602;
16'd13093 : result1 = 181615;
16'd13094 : result1 = 180602;
16'd13095 : result1 = 179561;
16'd13096 : result1 = 178491;
16'd13097 : result1 = 177391;
16'd13098 : result1 = 176258;
16'd13099 : result1 = 175091;
16'd13100 : result1 = 173886;
16'd13101 : result1 = 172642;
16'd13102 : result1 = 171354;
16'd13103 : result1 = 170018;
16'd13104 : result1 = 168631;
16'd13105 : result1 = 167186;
16'd13106 : result1 = 165677;
16'd13312 : result1 = 200628;
16'd13313 : result1 = 200584;
16'd13314 : result1 = 200497;
16'd13315 : result1 = 200371;
16'd13316 : result1 = 200206;
16'd13317 : result1 = 200005;
16'd13318 : result1 = 199770;
16'd13319 : result1 = 199502;
16'd13320 : result1 = 199203;
16'd13321 : result1 = 198873;
16'd13322 : result1 = 198515;
16'd13323 : result1 = 198129;
16'd13324 : result1 = 197716;
16'd13325 : result1 = 197278;
16'd13326 : result1 = 196814;
16'd13327 : result1 = 196327;
16'd13328 : result1 = 195816;
16'd13329 : result1 = 195281;
16'd13330 : result1 = 194725;
16'd13331 : result1 = 194146;
16'd13332 : result1 = 193546;
16'd13333 : result1 = 192925;
16'd13334 : result1 = 192283;
16'd13335 : result1 = 191619;
16'd13336 : result1 = 190935;
16'd13337 : result1 = 190231;
16'd13338 : result1 = 189505;
16'd13339 : result1 = 188759;
16'd13340 : result1 = 187992;
16'd13341 : result1 = 187204;
16'd13342 : result1 = 186394;
16'd13343 : result1 = 185563;
16'd13344 : result1 = 184709;
16'd13345 : result1 = 183832;
16'd13346 : result1 = 182932;
16'd13347 : result1 = 182008;
16'd13348 : result1 = 181059;
16'd13349 : result1 = 180083;
16'd13350 : result1 = 179081;
16'd13351 : result1 = 178049;
16'd13352 : result1 = 176988;
16'd13353 : result1 = 175895;
16'd13354 : result1 = 174769;
16'd13355 : result1 = 173607;
16'd13356 : result1 = 172406;
16'd13357 : result1 = 171163;
16'd13358 : result1 = 169875;
16'd13359 : result1 = 168539;
16'd13360 : result1 = 167147;
16'd13361 : result1 = 165696;
16'd13362 : result1 = 164177;
16'd13568 : result1 = 198082;
16'd13569 : result1 = 198081;
16'd13570 : result1 = 198037;
16'd13571 : result1 = 197953;
16'd13572 : result1 = 197829;
16'd13573 : result1 = 197669;
16'd13574 : result1 = 197474;
16'd13575 : result1 = 197244;
16'd13576 : result1 = 196983;
16'd13577 : result1 = 196690;
16'd13578 : result1 = 196367;
16'd13579 : result1 = 196016;
16'd13580 : result1 = 195637;
16'd13581 : result1 = 195231;
16'd13582 : result1 = 194799;
16'd13583 : result1 = 194342;
16'd13584 : result1 = 193860;
16'd13585 : result1 = 193355;
16'd13586 : result1 = 192826;
16'd13587 : result1 = 192274;
16'd13588 : result1 = 191700;
16'd13589 : result1 = 191103;
16'd13590 : result1 = 190485;
16'd13591 : result1 = 189845;
16'd13592 : result1 = 189183;
16'd13593 : result1 = 188500;
16'd13594 : result1 = 187795;
16'd13595 : result1 = 187068;
16'd13596 : result1 = 186320;
16'd13597 : result1 = 185550;
16'd13598 : result1 = 184757;
16'd13599 : result1 = 183942;
16'd13600 : result1 = 183103;
16'd13601 : result1 = 182241;
16'd13602 : result1 = 181355;
16'd13603 : result1 = 180443;
16'd13604 : result1 = 179506;
16'd13605 : result1 = 178541;
16'd13606 : result1 = 177548;
16'd13607 : result1 = 176526;
16'd13608 : result1 = 175472;
16'd13609 : result1 = 174386;
16'd13610 : result1 = 173265;
16'd13611 : result1 = 172107;
16'd13612 : result1 = 170908;
16'd13613 : result1 = 169667;
16'd13614 : result1 = 168378;
16'd13615 : result1 = 167038;
16'd13616 : result1 = 165642;
16'd13617 : result1 = 164182;
16'd13618 : result1 = 162652;
16'd13824 : result1 = 195591;
16'd13825 : result1 = 195629;
16'd13826 : result1 = 195624;
16'd13827 : result1 = 195578;
16'd13828 : result1 = 195492;
16'd13829 : result1 = 195369;
16'd13830 : result1 = 195210;
16'd13831 : result1 = 195017;
16'd13832 : result1 = 194790;
16'd13833 : result1 = 194531;
16'd13834 : result1 = 194242;
16'd13835 : result1 = 193923;
16'd13836 : result1 = 193575;
16'd13837 : result1 = 193200;
16'd13838 : result1 = 192798;
16'd13839 : result1 = 192369;
16'd13840 : result1 = 191916;
16'd13841 : result1 = 191437;
16'd13842 : result1 = 190935;
16'd13843 : result1 = 190408;
16'd13844 : result1 = 189859;
16'd13845 : result1 = 189286;
16'd13846 : result1 = 188690;
16'd13847 : result1 = 188072;
16'd13848 : result1 = 187431;
16'd13849 : result1 = 186768;
16'd13850 : result1 = 186083;
16'd13851 : result1 = 185375;
16'd13852 : result1 = 184645;
16'd13853 : result1 = 183891;
16'd13854 : result1 = 183115;
16'd13855 : result1 = 182315;
16'd13856 : result1 = 181491;
16'd13857 : result1 = 180643;
16'd13858 : result1 = 179769;
16'd13859 : result1 = 178869;
16'd13860 : result1 = 177943;
16'd13861 : result1 = 176988;
16'd13862 : result1 = 176004;
16'd13863 : result1 = 174990;
16'd13864 : result1 = 173944;
16'd13865 : result1 = 172863;
16'd13866 : result1 = 171746;
16'd13867 : result1 = 170591;
16'd13868 : result1 = 169394;
16'd13869 : result1 = 168152;
16'd13870 : result1 = 166861;
16'd13871 : result1 = 165517;
16'd13872 : result1 = 164113;
16'd13873 : result1 = 162643;
16'd13874 : result1 = 161099;
16'd14080 : result1 = 193153;
16'd14081 : result1 = 193226;
16'd14082 : result1 = 193256;
16'd14083 : result1 = 193245;
16'd14084 : result1 = 193194;
16'd14085 : result1 = 193105;
16'd14086 : result1 = 192979;
16'd14087 : result1 = 192818;
16'd14088 : result1 = 192624;
16'd14089 : result1 = 192397;
16'd14090 : result1 = 192138;
16'd14091 : result1 = 191849;
16'd14092 : result1 = 191531;
16'd14093 : result1 = 191185;
16'd14094 : result1 = 190810;
16'd14095 : result1 = 190409;
16'd14096 : result1 = 189982;
16'd14097 : result1 = 189529;
16'd14098 : result1 = 189052;
16'd14099 : result1 = 188549;
16'd14100 : result1 = 188023;
16'd14101 : result1 = 187472;
16'd14102 : result1 = 186898;
16'd14103 : result1 = 186301;
16'd14104 : result1 = 185680;
16'd14105 : result1 = 185037;
16'd14106 : result1 = 184370;
16'd14107 : result1 = 183680;
16'd14108 : result1 = 182966;
16'd14109 : result1 = 182229;
16'd14110 : result1 = 181468;
16'd14111 : result1 = 180683;
16'd14112 : result1 = 179872;
16'd14113 : result1 = 179037;
16'd14114 : result1 = 178175;
16'd14115 : result1 = 177287;
16'd14116 : result1 = 176370;
16'd14117 : result1 = 175425;
16'd14118 : result1 = 174449;
16'd14119 : result1 = 173442;
16'd14120 : result1 = 172401;
16'd14121 : result1 = 171326;
16'd14122 : result1 = 170212;
16'd14123 : result1 = 169059;
16'd14124 : result1 = 167862;
16'd14125 : result1 = 166618;
16'd14126 : result1 = 165324;
16'd14127 : result1 = 163973;
16'd14128 : result1 = 162560;
16'd14129 : result1 = 161078;
16'd14130 : result1 = 159516;
16'd14336 : result1 = 190765;
16'd14337 : result1 = 190870;
16'd14338 : result1 = 190932;
16'd14339 : result1 = 190952;
16'd14340 : result1 = 190932;
16'd14341 : result1 = 190874;
16'd14342 : result1 = 190779;
16'd14343 : result1 = 190649;
16'd14344 : result1 = 190484;
16'd14345 : result1 = 190286;
16'd14346 : result1 = 190056;
16'd14347 : result1 = 189796;
16'd14348 : result1 = 189505;
16'd14349 : result1 = 189185;
16'd14350 : result1 = 188837;
16'd14351 : result1 = 188462;
16'd14352 : result1 = 188059;
16'd14353 : result1 = 187631;
16'd14354 : result1 = 187176;
16'd14355 : result1 = 186696;
16'd14356 : result1 = 186192;
16'd14357 : result1 = 185663;
16'd14358 : result1 = 185109;
16'd14359 : result1 = 184532;
16'd14360 : result1 = 183930;
16'd14361 : result1 = 183305;
16'd14362 : result1 = 182655;
16'd14363 : result1 = 181982;
16'd14364 : result1 = 181285;
16'd14365 : result1 = 180563;
16'd14366 : result1 = 179816;
16'd14367 : result1 = 179044;
16'd14368 : result1 = 178247;
16'd14369 : result1 = 177424;
16'd14370 : result1 = 176573;
16'd14371 : result1 = 175695;
16'd14372 : result1 = 174788;
16'd14373 : result1 = 173851;
16'd14374 : result1 = 172882;
16'd14375 : result1 = 171881;
16'd14376 : result1 = 170846;
16'd14377 : result1 = 169773;
16'd14378 : result1 = 168662;
16'd14379 : result1 = 167509;
16'd14380 : result1 = 166311;
16'd14381 : result1 = 165065;
16'd14382 : result1 = 163765;
16'd14383 : result1 = 162406;
16'd14384 : result1 = 160982;
16'd14385 : result1 = 159484;
16'd14386 : result1 = 157903;
16'd14592 : result1 = 188425;
16'd14593 : result1 = 188559;
16'd14594 : result1 = 188649;
16'd14595 : result1 = 188697;
16'd14596 : result1 = 188706;
16'd14597 : result1 = 188677;
16'd14598 : result1 = 188610;
16'd14599 : result1 = 188507;
16'd14600 : result1 = 188370;
16'd14601 : result1 = 188199;
16'd14602 : result1 = 187996;
16'd14603 : result1 = 187761;
16'd14604 : result1 = 187496;
16'd14605 : result1 = 187201;
16'd14606 : result1 = 186878;
16'd14607 : result1 = 186526;
16'd14608 : result1 = 186147;
16'd14609 : result1 = 185741;
16'd14610 : result1 = 185309;
16'd14611 : result1 = 184850;
16'd14612 : result1 = 184366;
16'd14613 : result1 = 183857;
16'd14614 : result1 = 183323;
16'd14615 : result1 = 182764;
16'd14616 : result1 = 182181;
16'd14617 : result1 = 181573;
16'd14618 : result1 = 180940;
16'd14619 : result1 = 180282;
16'd14620 : result1 = 179600;
16'd14621 : result1 = 178892;
16'd14622 : result1 = 178159;
16'd14623 : result1 = 177401;
16'd14624 : result1 = 176615;
16'd14625 : result1 = 175803;
16'd14626 : result1 = 174963;
16'd14627 : result1 = 174094;
16'd14628 : result1 = 173195;
16'd14629 : result1 = 172265;
16'd14630 : result1 = 171303;
16'd14631 : result1 = 170307;
16'd14632 : result1 = 169276;
16'd14633 : result1 = 168206;
16'd14634 : result1 = 167096;
16'd14635 : result1 = 165942;
16'd14636 : result1 = 164742;
16'd14637 : result1 = 163490;
16'd14638 : result1 = 162183;
16'd14639 : result1 = 160814;
16'd14640 : result1 = 159376;
16'd14641 : result1 = 157861;
16'd14642 : result1 = 156256;
16'd14848 : result1 = 186131;
16'd14849 : result1 = 186290;
16'd14850 : result1 = 186405;
16'd14851 : result1 = 186480;
16'd14852 : result1 = 186514;
16'd14853 : result1 = 186510;
16'd14854 : result1 = 186469;
16'd14855 : result1 = 186392;
16'd14856 : result1 = 186280;
16'd14857 : result1 = 186134;
16'd14858 : result1 = 185956;
16'd14859 : result1 = 185745;
16'd14860 : result1 = 185504;
16'd14861 : result1 = 185233;
16'd14862 : result1 = 184932;
16'd14863 : result1 = 184603;
16'd14864 : result1 = 184245;
16'd14865 : result1 = 183860;
16'd14866 : result1 = 183449;
16'd14867 : result1 = 183011;
16'd14868 : result1 = 182546;
16'd14869 : result1 = 182056;
16'd14870 : result1 = 181540;
16'd14871 : result1 = 180999;
16'd14872 : result1 = 180432;
16'd14873 : result1 = 179840;
16'd14874 : result1 = 179223;
16'd14875 : result1 = 178580;
16'd14876 : result1 = 177912;
16'd14877 : result1 = 177218;
16'd14878 : result1 = 176498;
16'd14879 : result1 = 175751;
16'd14880 : result1 = 174976;
16'd14881 : result1 = 174174;
16'd14882 : result1 = 173343;
16'd14883 : result1 = 172483;
16'd14884 : result1 = 171592;
16'd14885 : result1 = 170668;
16'd14886 : result1 = 169712;
16'd14887 : result1 = 168720;
16'd14888 : result1 = 167691;
16'd14889 : result1 = 166623;
16'd14890 : result1 = 165512;
16'd14891 : result1 = 164357;
16'd14892 : result1 = 163152;
16'd14893 : result1 = 161894;
16'd14894 : result1 = 160577;
16'd14895 : result1 = 159196;
16'd14896 : result1 = 157742;
16'd14897 : result1 = 156205;
16'd14898 : result1 = 154574;
16'd15104 : result1 = 183880;
16'd15105 : result1 = 184061;
16'd15106 : result1 = 184200;
16'd15107 : result1 = 184297;
16'd15108 : result1 = 184355;
16'd15109 : result1 = 184375;
16'd15110 : result1 = 184357;
16'd15111 : result1 = 184303;
16'd15112 : result1 = 184214;
16'd15113 : result1 = 184091;
16'd15114 : result1 = 183935;
16'd15115 : result1 = 183747;
16'd15116 : result1 = 183528;
16'd15117 : result1 = 183279;
16'd15118 : result1 = 182999;
16'd15119 : result1 = 182691;
16'd15120 : result1 = 182354;
16'd15121 : result1 = 181989;
16'd15122 : result1 = 181596;
16'd15123 : result1 = 181177;
16'd15124 : result1 = 180731;
16'd15125 : result1 = 180258;
16'd15126 : result1 = 179760;
16'd15127 : result1 = 179235;
16'd15128 : result1 = 178684;
16'd15129 : result1 = 178107;
16'd15130 : result1 = 177505;
16'd15131 : result1 = 176876;
16'd15132 : result1 = 176221;
16'd15133 : result1 = 175540;
16'd15134 : result1 = 174831;
16'd15135 : result1 = 174095;
16'd15136 : result1 = 173331;
16'd15137 : result1 = 172538;
16'd15138 : result1 = 171715;
16'd15139 : result1 = 170862;
16'd15140 : result1 = 169978;
16'd15141 : result1 = 169060;
16'd15142 : result1 = 168107;
16'd15143 : result1 = 167119;
16'd15144 : result1 = 166091;
16'd15145 : result1 = 165023;
16'd15146 : result1 = 163911;
16'd15147 : result1 = 162751;
16'd15148 : result1 = 161541;
16'd15149 : result1 = 160275;
16'd15150 : result1 = 158947;
16'd15151 : result1 = 157550;
16'd15152 : result1 = 156076;
16'd15153 : result1 = 154515;
16'd15154 : result1 = 152851;
16'd15360 : result1 = 181670;
16'd15361 : result1 = 181871;
16'd15362 : result1 = 182030;
16'd15363 : result1 = 182148;
16'd15364 : result1 = 182227;
16'd15365 : result1 = 182268;
16'd15366 : result1 = 182271;
16'd15367 : result1 = 182239;
16'd15368 : result1 = 182171;
16'd15369 : result1 = 182069;
16'd15370 : result1 = 181934;
16'd15371 : result1 = 181767;
16'd15372 : result1 = 181568;
16'd15373 : result1 = 181339;
16'd15374 : result1 = 181079;
16'd15375 : result1 = 180790;
16'd15376 : result1 = 180472;
16'd15377 : result1 = 180126;
16'd15378 : result1 = 179752;
16'd15379 : result1 = 179350;
16'd15380 : result1 = 178921;
16'd15381 : result1 = 178465;
16'd15382 : result1 = 177982;
16'd15383 : result1 = 177472;
16'd15384 : result1 = 176937;
16'd15385 : result1 = 176374;
16'd15386 : result1 = 175785;
16'd15387 : result1 = 175169;
16'd15388 : result1 = 174527;
16'd15389 : result1 = 173856;
16'd15390 : result1 = 173159;
16'd15391 : result1 = 172433;
16'd15392 : result1 = 171678;
16'd15393 : result1 = 170893;
16'd15394 : result1 = 170078;
16'd15395 : result1 = 169232;
16'd15396 : result1 = 168352;
16'd15397 : result1 = 167439;
16'd15398 : result1 = 166489;
16'd15399 : result1 = 165502;
16'd15400 : result1 = 164475;
16'd15401 : result1 = 163406;
16'd15402 : result1 = 162290;
16'd15403 : result1 = 161126;
16'd15404 : result1 = 159907;
16'd15405 : result1 = 158631;
16'd15406 : result1 = 157289;
16'd15407 : result1 = 155874;
16'd15408 : result1 = 154378;
16'd15409 : result1 = 152787;
16'd15410 : result1 = 151086;
16'd15616 : result1 = 179498;
16'd15617 : result1 = 179717;
16'd15618 : result1 = 179894;
16'd15619 : result1 = 180031;
16'd15620 : result1 = 180129;
16'd15621 : result1 = 180189;
16'd15622 : result1 = 180212;
16'd15623 : result1 = 180198;
16'd15624 : result1 = 180150;
16'd15625 : result1 = 180068;
16'd15626 : result1 = 179952;
16'd15627 : result1 = 179804;
16'd15628 : result1 = 179624;
16'd15629 : result1 = 179413;
16'd15630 : result1 = 179172;
16'd15631 : result1 = 178901;
16'd15632 : result1 = 178600;
16'd15633 : result1 = 178271;
16'd15634 : result1 = 177914;
16'd15635 : result1 = 177528;
16'd15636 : result1 = 177115;
16'd15637 : result1 = 176674;
16'd15638 : result1 = 176206;
16'd15639 : result1 = 175711;
16'd15640 : result1 = 175189;
16'd15641 : result1 = 174640;
16'd15642 : result1 = 174064;
16'd15643 : result1 = 173460;
16'd15644 : result1 = 172828;
16'd15645 : result1 = 172169;
16'd15646 : result1 = 171481;
16'd15647 : result1 = 170764;
16'd15648 : result1 = 170017;
16'd15649 : result1 = 169240;
16'd15650 : result1 = 168431;
16'd15651 : result1 = 167590;
16'd15652 : result1 = 166715;
16'd15653 : result1 = 165805;
16'd15654 : result1 = 164857;
16'd15655 : result1 = 163871;
16'd15656 : result1 = 162842;
16'd15657 : result1 = 161770;
16'd15658 : result1 = 160650;
16'd15659 : result1 = 159478;
16'd15660 : result1 = 158250;
16'd15661 : result1 = 156960;
16'd15662 : result1 = 155602;
16'd15663 : result1 = 154166;
16'd15664 : result1 = 152642;
16'd15665 : result1 = 151017;
16'd15666 : result1 = 149272;
16'd15872 : result1 = 177363;
16'd15873 : result1 = 177597;
16'd15874 : result1 = 177791;
16'd15875 : result1 = 177944;
16'd15876 : result1 = 178059;
16'd15877 : result1 = 178136;
16'd15878 : result1 = 178176;
16'd15879 : result1 = 178181;
16'd15880 : result1 = 178150;
16'd15881 : result1 = 178085;
16'd15882 : result1 = 177987;
16'd15883 : result1 = 177857;
16'd15884 : result1 = 177694;
16'd15885 : result1 = 177500;
16'd15886 : result1 = 177276;
16'd15887 : result1 = 177021;
16'd15888 : result1 = 176737;
16'd15889 : result1 = 176424;
16'd15890 : result1 = 176082;
16'd15891 : result1 = 175712;
16'd15892 : result1 = 175313;
16'd15893 : result1 = 174887;
16'd15894 : result1 = 174433;
16'd15895 : result1 = 173951;
16'd15896 : result1 = 173442;
16'd15897 : result1 = 172905;
16'd15898 : result1 = 172340;
16'd15899 : result1 = 171747;
16'd15900 : result1 = 171126;
16'd15901 : result1 = 170476;
16'd15902 : result1 = 169797;
16'd15903 : result1 = 169088;
16'd15904 : result1 = 168348;
16'd15905 : result1 = 167577;
16'd15906 : result1 = 166774;
16'd15907 : result1 = 165937;
16'd15908 : result1 = 165065;
16'd15909 : result1 = 164157;
16'd15910 : result1 = 163210;
16'd15911 : result1 = 162223;
16'd15912 : result1 = 161192;
16'd15913 : result1 = 160115;
16'd15914 : result1 = 158988;
16'd15915 : result1 = 157807;
16'd15916 : result1 = 156567;
16'd15917 : result1 = 155261;
16'd15918 : result1 = 153883;
16'd15919 : result1 = 152422;
16'd15920 : result1 = 150867;
16'd15921 : result1 = 149201;
16'd15922 : result1 = 147405;
16'd16128 : result1 = 175262;
16'd16129 : result1 = 175510;
16'd16130 : result1 = 175718;
16'd16131 : result1 = 175886;
16'd16132 : result1 = 176016;
16'd16133 : result1 = 176108;
16'd16134 : result1 = 176164;
16'd16135 : result1 = 176185;
16'd16136 : result1 = 176170;
16'd16137 : result1 = 176121;
16'd16138 : result1 = 176039;
16'd16139 : result1 = 175925;
16'd16140 : result1 = 175778;
16'd16141 : result1 = 175600;
16'd16142 : result1 = 175391;
16'd16143 : result1 = 175152;
16'd16144 : result1 = 174883;
16'd16145 : result1 = 174584;
16'd16146 : result1 = 174257;
16'd16147 : result1 = 173901;
16'd16148 : result1 = 173516;
16'd16149 : result1 = 173103;
16'd16150 : result1 = 172661;
16'd16151 : result1 = 172192;
16'd16152 : result1 = 171694;
16'd16153 : result1 = 171168;
16'd16154 : result1 = 170614;
16'd16155 : result1 = 170031;
16'd16156 : result1 = 169419;
16'd16157 : result1 = 168777;
16'd16158 : result1 = 168106;
16'd16159 : result1 = 167404;
16'd16160 : result1 = 166671;
16'd16161 : result1 = 165905;
16'd16162 : result1 = 165106;
16'd16163 : result1 = 164272;
16'd16164 : result1 = 163402;
16'd16165 : result1 = 162495;
16'd16166 : result1 = 161547;
16'd16167 : result1 = 160557;
16'd16168 : result1 = 159522;
16'd16169 : result1 = 158439;
16'd16170 : result1 = 157303;
16'd16171 : result1 = 156111;
16'd16172 : result1 = 154856;
16'd16173 : result1 = 153532;
16'd16174 : result1 = 152130;
16'd16175 : result1 = 150640;
16'd16176 : result1 = 149047;
16'd16177 : result1 = 147335;
16'd16178 : result1 = 145477;
16'd16384 : result1 = 173193;
16'd16385 : result1 = 173453;
16'd16386 : result1 = 173673;
16'd16387 : result1 = 173855;
16'd16388 : result1 = 173998;
16'd16389 : result1 = 174104;
16'd16390 : result1 = 174175;
16'd16391 : result1 = 174209;
16'd16392 : result1 = 174209;
16'd16393 : result1 = 174175;
16'd16394 : result1 = 174108;
16'd16395 : result1 = 174007;
16'd16396 : result1 = 173875;
16'd16397 : result1 = 173712;
16'd16398 : result1 = 173517;
16'd16399 : result1 = 173292;
16'd16400 : result1 = 173037;
16'd16401 : result1 = 172752;
16'd16402 : result1 = 172437;
16'd16403 : result1 = 172094;
16'd16404 : result1 = 171722;
16'd16405 : result1 = 171320;
16'd16406 : result1 = 170891;
16'd16407 : result1 = 170432;
16'd16408 : result1 = 169945;
16'd16409 : result1 = 169429;
16'd16410 : result1 = 168885;
16'd16411 : result1 = 168310;
16'd16412 : result1 = 167707;
16'd16413 : result1 = 167073;
16'd16414 : result1 = 166408;
16'd16415 : result1 = 165712;
16'd16416 : result1 = 164984;
16'd16417 : result1 = 164222;
16'd16418 : result1 = 163426;
16'd16419 : result1 = 162595;
16'd16420 : result1 = 161725;
16'd16421 : result1 = 160817;
16'd16422 : result1 = 159867;
16'd16423 : result1 = 158873;
16'd16424 : result1 = 157832;
16'd16425 : result1 = 156741;
16'd16426 : result1 = 155594;
16'd16427 : result1 = 154388;
16'd16428 : result1 = 153115;
16'd16429 : result1 = 151769;
16'd16430 : result1 = 150339;
16'd16431 : result1 = 148814;
16'd16432 : result1 = 147178;
16'd16433 : result1 = 145410;
16'd16434 : result1 = 143480;
16'd16640 : result1 = 171154;
16'd16641 : result1 = 171425;
16'd16642 : result1 = 171656;
16'd16643 : result1 = 171849;
16'd16644 : result1 = 172004;
16'd16645 : result1 = 172123;
16'd16646 : result1 = 172206;
16'd16647 : result1 = 172253;
16'd16648 : result1 = 172266;
16'd16649 : result1 = 172245;
16'd16650 : result1 = 172191;
16'd16651 : result1 = 172104;
16'd16652 : result1 = 171985;
16'd16653 : result1 = 171834;
16'd16654 : result1 = 171653;
16'd16655 : result1 = 171440;
16'd16656 : result1 = 171198;
16'd16657 : result1 = 170925;
16'd16658 : result1 = 170623;
16'd16659 : result1 = 170291;
16'd16660 : result1 = 169930;
16'd16661 : result1 = 169540;
16'd16662 : result1 = 169121;
16'd16663 : result1 = 168673;
16'd16664 : result1 = 168195;
16'd16665 : result1 = 167688;
16'd16666 : result1 = 167152;
16'd16667 : result1 = 166586;
16'd16668 : result1 = 165989;
16'd16669 : result1 = 165362;
16'd16670 : result1 = 164703;
16'd16671 : result1 = 164011;
16'd16672 : result1 = 163287;
16'd16673 : result1 = 162528;
16'd16674 : result1 = 161734;
16'd16675 : result1 = 160903;
16'd16676 : result1 = 160033;
16'd16677 : result1 = 159123;
16'd16678 : result1 = 158169;
16'd16679 : result1 = 157169;
16'd16680 : result1 = 156120;
16'd16681 : result1 = 155018;
16'd16682 : result1 = 153858;
16'd16683 : result1 = 152635;
16'd16684 : result1 = 151342;
16'd16685 : result1 = 149969;
16'd16686 : result1 = 148507;
16'd16687 : result1 = 146941;
16'd16688 : result1 = 145254;
16'd16689 : result1 = 143419;
16'd16690 : result1 = 141401;
16'd16896 : result1 = 169144;
16'd16897 : result1 = 169423;
16'd16898 : result1 = 169664;
16'd16899 : result1 = 169867;
16'd16900 : result1 = 170033;
16'd16901 : result1 = 170162;
16'd16902 : result1 = 170256;
16'd16903 : result1 = 170315;
16'd16904 : result1 = 170340;
16'd16905 : result1 = 170330;
16'd16906 : result1 = 170288;
16'd16907 : result1 = 170213;
16'd16908 : result1 = 170106;
16'd16909 : result1 = 169967;
16'd16910 : result1 = 169798;
16'd16911 : result1 = 169597;
16'd16912 : result1 = 169366;
16'd16913 : result1 = 169104;
16'd16914 : result1 = 168813;
16'd16915 : result1 = 168492;
16'd16916 : result1 = 168141;
16'd16917 : result1 = 167761;
16'd16918 : result1 = 167351;
16'd16919 : result1 = 166912;
16'd16920 : result1 = 166443;
16'd16921 : result1 = 165944;
16'd16922 : result1 = 165415;
16'd16923 : result1 = 164856;
16'd16924 : result1 = 164265;
16'd16925 : result1 = 163643;
16'd16926 : result1 = 162989;
16'd16927 : result1 = 162301;
16'd16928 : result1 = 161580;
16'd16929 : result1 = 160823;
16'd16930 : result1 = 160029;
16'd16931 : result1 = 159197;
16'd16932 : result1 = 158325;
16'd16933 : result1 = 157411;
16'd16934 : result1 = 156451;
16'd16935 : result1 = 155444;
16'd16936 : result1 = 154385;
16'd16937 : result1 = 153270;
16'd16938 : result1 = 152094;
16'd16939 : result1 = 150851;
16'd16940 : result1 = 149532;
16'd16941 : result1 = 148129;
16'd16942 : result1 = 146629;
16'd16943 : result1 = 145015;
16'd16944 : result1 = 143266;
16'd16945 : result1 = 141351;
16'd16946 : result1 = 139226;
16'd17152 : result1 = 167160;
16'd17153 : result1 = 167447;
16'd17154 : result1 = 167695;
16'd17155 : result1 = 167907;
16'd17156 : result1 = 168082;
16'd17157 : result1 = 168221;
16'd17158 : result1 = 168325;
16'd17159 : result1 = 168394;
16'd17160 : result1 = 168429;
16'd17161 : result1 = 168430;
16'd17162 : result1 = 168399;
16'd17163 : result1 = 168334;
16'd17164 : result1 = 168238;
16'd17165 : result1 = 168110;
16'd17166 : result1 = 167951;
16'd17167 : result1 = 167760;
16'd17168 : result1 = 167539;
16'd17169 : result1 = 167288;
16'd17170 : result1 = 167007;
16'd17171 : result1 = 166695;
16'd17172 : result1 = 166354;
16'd17173 : result1 = 165982;
16'd17174 : result1 = 165581;
16'd17175 : result1 = 165150;
16'd17176 : result1 = 164688;
16'd17177 : result1 = 164196;
16'd17178 : result1 = 163674;
16'd17179 : result1 = 163120;
16'd17180 : result1 = 162534;
16'd17181 : result1 = 161917;
16'd17182 : result1 = 161266;
16'd17183 : result1 = 160581;
16'd17184 : result1 = 159860;
16'd17185 : result1 = 159104;
16'd17186 : result1 = 158309;
16'd17187 : result1 = 157475;
16'd17188 : result1 = 156599;
16'd17189 : result1 = 155679;
16'd17190 : result1 = 154712;
16'd17191 : result1 = 153695;
16'd17192 : result1 = 152624;
16'd17193 : result1 = 151493;
16'd17194 : result1 = 150298;
16'd17195 : result1 = 149031;
16'd17196 : result1 = 147683;
16'd17197 : result1 = 146244;
16'd17198 : result1 = 144698;
16'd17199 : result1 = 143027;
16'd17200 : result1 = 141205;
16'd17201 : result1 = 139193;
16'd17202 : result1 = 136934;
16'd17408 : result1 = 165200;
16'd17409 : result1 = 165493;
16'd17410 : result1 = 165749;
16'd17411 : result1 = 165968;
16'd17412 : result1 = 166151;
16'd17413 : result1 = 166298;
16'd17414 : result1 = 166411;
16'd17415 : result1 = 166489;
16'd17416 : result1 = 166533;
16'd17417 : result1 = 166544;
16'd17418 : result1 = 166521;
16'd17419 : result1 = 166467;
16'd17420 : result1 = 166380;
16'd17421 : result1 = 166261;
16'd17422 : result1 = 166111;
16'd17423 : result1 = 165930;
16'd17424 : result1 = 165719;
16'd17425 : result1 = 165476;
16'd17426 : result1 = 165204;
16'd17427 : result1 = 164901;
16'd17428 : result1 = 164567;
16'd17429 : result1 = 164204;
16'd17430 : result1 = 163810;
16'd17431 : result1 = 163385;
16'd17432 : result1 = 162930;
16'd17433 : result1 = 162444;
16'd17434 : result1 = 161927;
16'd17435 : result1 = 161378;
16'd17436 : result1 = 160796;
16'd17437 : result1 = 160181;
16'd17438 : result1 = 159532;
16'd17439 : result1 = 158848;
16'd17440 : result1 = 158128;
16'd17441 : result1 = 157371;
16'd17442 : result1 = 156574;
16'd17443 : result1 = 155736;
16'd17444 : result1 = 154854;
16'd17445 : result1 = 153927;
16'd17446 : result1 = 152950;
16'd17447 : result1 = 151921;
16'd17448 : result1 = 150834;
16'd17449 : result1 = 149685;
16'd17450 : result1 = 148467;
16'd17451 : result1 = 147172;
16'd17452 : result1 = 145790;
16'd17453 : result1 = 144308;
16'd17454 : result1 = 142709;
16'd17455 : result1 = 140970;
16'd17456 : result1 = 139058;
16'd17457 : result1 = 136926;
16'd17458 : result1 = 134497;
16'd17664 : result1 = 163264;
16'd17665 : result1 = 163562;
16'd17666 : result1 = 163823;
16'd17667 : result1 = 164048;
16'd17668 : result1 = 164238;
16'd17669 : result1 = 164392;
16'd17670 : result1 = 164512;
16'd17671 : result1 = 164598;
16'd17672 : result1 = 164650;
16'd17673 : result1 = 164669;
16'd17674 : result1 = 164655;
16'd17675 : result1 = 164609;
16'd17676 : result1 = 164530;
16'd17677 : result1 = 164420;
16'd17678 : result1 = 164279;
16'd17679 : result1 = 164106;
16'd17680 : result1 = 163902;
16'd17681 : result1 = 163668;
16'd17682 : result1 = 163403;
16'd17683 : result1 = 163107;
16'd17684 : result1 = 162781;
16'd17685 : result1 = 162424;
16'd17686 : result1 = 162036;
16'd17687 : result1 = 161618;
16'd17688 : result1 = 161168;
16'd17689 : result1 = 160687;
16'd17690 : result1 = 160173;
16'd17691 : result1 = 159628;
16'd17692 : result1 = 159049;
16'd17693 : result1 = 158436;
16'd17694 : result1 = 157788;
16'd17695 : result1 = 157104;
16'd17696 : result1 = 156382;
16'd17697 : result1 = 155622;
16'd17698 : result1 = 154821;
16'd17699 : result1 = 153978;
16'd17700 : result1 = 153089;
16'd17701 : result1 = 152152;
16'd17702 : result1 = 151163;
16'd17703 : result1 = 150119;
16'd17704 : result1 = 149015;
16'd17705 : result1 = 147843;
16'd17706 : result1 = 146598;
16'd17707 : result1 = 145270;
16'd17708 : result1 = 143847;
16'd17709 : result1 = 142314;
16'd17710 : result1 = 140651;
16'd17711 : result1 = 138830;
16'd17712 : result1 = 136809;
16'd17713 : result1 = 134525;
16'd17714 : result1 = 131868;
16'd17920 : result1 = 161348;
16'd17921 : result1 = 161650;
16'd17922 : result1 = 161916;
16'd17923 : result1 = 162146;
16'd17924 : result1 = 162342;
16'd17925 : result1 = 162502;
16'd17926 : result1 = 162628;
16'd17927 : result1 = 162721;
16'd17928 : result1 = 162780;
16'd17929 : result1 = 162806;
16'd17930 : result1 = 162799;
16'd17931 : result1 = 162760;
16'd17932 : result1 = 162689;
16'd17933 : result1 = 162586;
16'd17934 : result1 = 162452;
16'd17935 : result1 = 162286;
16'd17936 : result1 = 162090;
16'd17937 : result1 = 161862;
16'd17938 : result1 = 161604;
16'd17939 : result1 = 161314;
16'd17940 : result1 = 160994;
16'd17941 : result1 = 160643;
16'd17942 : result1 = 160260;
16'd17943 : result1 = 159846;
16'd17944 : result1 = 159401;
16'd17945 : result1 = 158923;
16'd17946 : result1 = 158413;
16'd17947 : result1 = 157869;
16'd17948 : result1 = 157292;
16'd17949 : result1 = 156679;
16'd17950 : result1 = 156031;
16'd17951 : result1 = 155345;
16'd17952 : result1 = 154621;
16'd17953 : result1 = 153857;
16'd17954 : result1 = 153050;
16'd17955 : result1 = 152199;
16'd17956 : result1 = 151301;
16'd17957 : result1 = 150352;
16'd17958 : result1 = 149349;
16'd17959 : result1 = 148287;
16'd17960 : result1 = 147161;
16'd17961 : result1 = 145963;
16'd17962 : result1 = 144686;
16'd17963 : result1 = 143319;
16'd17964 : result1 = 141847;
16'd17965 : result1 = 140254;
16'd17966 : result1 = 138514;
16'd17967 : result1 = 136592;
16'd17968 : result1 = 134434;
16'd17969 : result1 = 131951;
16'd17970 : result1 = 128978;
16'd19758 : result1 = 118000;
endcase;

case(xy)

		16'd0 : result2 = 150955;
		16'd1 : result2 = 150776;
		16'd2 : result2 = 150567;
		16'd3 : result2 = 150330;
		16'd4 : result2 = 150073;
		16'd5 : result2 = 149798;
		16'd6 : result2 = 149511;
		16'd7 : result2 = 149216;
		16'd8 : result2 = 148915;
		16'd9 : result2 = 148612;
		16'd10 : result2 = 148310;
		16'd11 : result2 = 148012;
		16'd12 : result2 = 147721;
		16'd13 : result2 = 147437;
		16'd14 : result2 = 147165;
		16'd15 : result2 = 146904;
		16'd16 : result2 = 146658;
		16'd17 : result2 = 146426;
		16'd18 : result2 = 146212;
		16'd19 : result2 = 146015;
		16'd20 : result2 = 145837;
		16'd21 : result2 = 145679;
		16'd22 : result2 = 145542;
		16'd23 : result2 = 145427;
		16'd24 : result2 = 145334;
		16'd25 : result2 = 145265;
		16'd26 : result2 = 145219;
		16'd27 : result2 = 145198;
		16'd28 : result2 = 145203;
		16'd29 : result2 = 145234;
		16'd30 : result2 = 145291;
		16'd31 : result2 = 145376;
		16'd32 : result2 = 145489;
		16'd33 : result2 = 145632;
		16'd34 : result2 = 145804;
		16'd35 : result2 = 146007;
		16'd36 : result2 = 146242;
		16'd37 : result2 = 146510;
		16'd38 : result2 = 146812;
		16'd39 : result2 = 147150;
		16'd40 : result2 = 147526;
		16'd41 : result2 = 147940;
		16'd42 : result2 = 148397;
		16'd43 : result2 = 148897;
		16'd44 : result2 = 149444;
		16'd45 : result2 = 150041;
		16'd46 : result2 = 150693;
		16'd47 : result2 = 151404;
		16'd48 : result2 = 152181;
		16'd49 : result2 = 153031;
		16'd50 : result2 = 153963;
		16'd256 : result2 = 149173;
		16'd257 : result2 = 149035;
		16'd258 : result2 = 148858;
		16'd259 : result2 = 148649;
		16'd260 : result2 = 148413;
		16'd261 : result2 = 148156;
		16'd262 : result2 = 147882;
		16'd263 : result2 = 147597;
		16'd264 : result2 = 147304;
		16'd265 : result2 = 147007;
		16'd266 : result2 = 146710;
		16'd267 : result2 = 146415;
		16'd268 : result2 = 146125;
		16'd269 : result2 = 145843;
		16'd270 : result2 = 145571;
		16'd271 : result2 = 145310;
		16'd272 : result2 = 145063;
		16'd273 : result2 = 144831;
		16'd274 : result2 = 144615;
		16'd275 : result2 = 144416;
		16'd276 : result2 = 144237;
		16'd277 : result2 = 144077;
		16'd278 : result2 = 143938;
		16'd279 : result2 = 143821;
		16'd280 : result2 = 143725;
		16'd281 : result2 = 143653;
		16'd282 : result2 = 143605;
		16'd283 : result2 = 143581;
		16'd284 : result2 = 143583;
		16'd285 : result2 = 143610;
		16'd286 : result2 = 143664;
		16'd287 : result2 = 143744;
		16'd288 : result2 = 143853;
		16'd289 : result2 = 143990;
		16'd290 : result2 = 144156;
		16'd291 : result2 = 144353;
		16'd292 : result2 = 144581;
		16'd293 : result2 = 144841;
		16'd294 : result2 = 145134;
		16'd295 : result2 = 145462;
		16'd296 : result2 = 145827;
		16'd297 : result2 = 146229;
		16'd298 : result2 = 146671;
		16'd299 : result2 = 147154;
		16'd300 : result2 = 147683;
		16'd301 : result2 = 148259;
		16'd302 : result2 = 148886;
		16'd303 : result2 = 149570;
		16'd304 : result2 = 150314;
		16'd305 : result2 = 151125;
		16'd306 : result2 = 152011;
		16'd512 : result2 = 147380;
		16'd513 : result2 = 147287;
		16'd514 : result2 = 147147;
		16'd515 : result2 = 146967;
		16'd516 : result2 = 146754;
		16'd517 : result2 = 146515;
		16'd518 : result2 = 146255;
		16'd519 : result2 = 145981;
		16'd520 : result2 = 145697;
		16'd521 : result2 = 145406;
		16'd522 : result2 = 145113;
		16'd523 : result2 = 144821;
		16'd524 : result2 = 144534;
		16'd525 : result2 = 144253;
		16'd526 : result2 = 143981;
		16'd527 : result2 = 143720;
		16'd528 : result2 = 143473;
		16'd529 : result2 = 143240;
		16'd530 : result2 = 143023;
		16'd531 : result2 = 142823;
		16'd532 : result2 = 142642;
		16'd533 : result2 = 142481;
		16'd534 : result2 = 142341;
		16'd535 : result2 = 142221;
		16'd536 : result2 = 142124;
		16'd537 : result2 = 142050;
		16'd538 : result2 = 142000;
		16'd539 : result2 = 141974;
		16'd540 : result2 = 141973;
		16'd541 : result2 = 141997;
		16'd542 : result2 = 142048;
		16'd543 : result2 = 142125;
		16'd544 : result2 = 142230;
		16'd545 : result2 = 142363;
		16'd546 : result2 = 142524;
		16'd547 : result2 = 142716;
		16'd548 : result2 = 142938;
		16'd549 : result2 = 143191;
		16'd550 : result2 = 143477;
		16'd551 : result2 = 143796;
		16'd552 : result2 = 144151;
		16'd553 : result2 = 144542;
		16'd554 : result2 = 144971;
		16'd555 : result2 = 145441;
		16'd556 : result2 = 145954;
		16'd557 : result2 = 146511;
		16'd558 : result2 = 147118;
		16'd559 : result2 = 147777;
		16'd560 : result2 = 148493;
		16'd561 : result2 = 149271;
		16'd562 : result2 = 150119;
		16'd768 : result2 = 145577;
		16'd769 : result2 = 145534;
		16'd770 : result2 = 145434;
		16'd771 : result2 = 145285;
		16'd772 : result2 = 145096;
		16'd773 : result2 = 144876;
		16'd774 : result2 = 144631;
		16'd775 : result2 = 144368;
		16'd776 : result2 = 144092;
		16'd777 : result2 = 143808;
		16'd778 : result2 = 143520;
		16'd779 : result2 = 143231;
		16'd780 : result2 = 142946;
		16'd781 : result2 = 142666;
		16'd782 : result2 = 142395;
		16'd783 : result2 = 142134;
		16'd784 : result2 = 141886;
		16'd785 : result2 = 141653;
		16'd786 : result2 = 141435;
		16'd787 : result2 = 141235;
		16'd788 : result2 = 141053;
		16'd789 : result2 = 140891;
		16'd790 : result2 = 140749;
		16'd791 : result2 = 140628;
		16'd792 : result2 = 140530;
		16'd793 : result2 = 140454;
		16'd794 : result2 = 140402;
		16'd795 : result2 = 140375;
		16'd796 : result2 = 140372;
		16'd797 : result2 = 140394;
		16'd798 : result2 = 140442;
		16'd799 : result2 = 140517;
		16'd800 : result2 = 140619;
		16'd801 : result2 = 140748;
		16'd802 : result2 = 140906;
		16'd803 : result2 = 141093;
		16'd804 : result2 = 141310;
		16'd805 : result2 = 141558;
		16'd806 : result2 = 141837;
		16'd807 : result2 = 142150;
		16'd808 : result2 = 142496;
		16'd809 : result2 = 142878;
		16'd810 : result2 = 143297;
		16'd811 : result2 = 143754;
		16'd812 : result2 = 144253;
		16'd813 : result2 = 144795;
		16'd814 : result2 = 145383;
		16'd815 : result2 = 146021;
		16'd816 : result2 = 146713;
		16'd817 : result2 = 147463;
		16'd818 : result2 = 148277;
		16'd1024 : result2 = 143767;
		16'd1025 : result2 = 143778;
		16'd1026 : result2 = 143720;
		16'd1027 : result2 = 143604;
		16'd1028 : result2 = 143441;
		16'd1029 : result2 = 143241;
		16'd1030 : result2 = 143011;
		16'd1031 : result2 = 142759;
		16'd1032 : result2 = 142492;
		16'd1033 : result2 = 142214;
		16'd1034 : result2 = 141930;
		16'd1035 : result2 = 141644;
		16'd1036 : result2 = 141361;
		16'd1037 : result2 = 141082;
		16'd1038 : result2 = 140812;
		16'd1039 : result2 = 140551;
		16'd1040 : result2 = 140303;
		16'd1041 : result2 = 140070;
		16'd1042 : result2 = 139851;
		16'd1043 : result2 = 139650;
		16'd1044 : result2 = 139468;
		16'd1045 : result2 = 139305;
		16'd1046 : result2 = 139162;
		16'd1047 : result2 = 139041;
		16'd1048 : result2 = 138941;
		16'd1049 : result2 = 138865;
		16'd1050 : result2 = 138812;
		16'd1051 : result2 = 138783;
		16'd1052 : result2 = 138778;
		16'd1053 : result2 = 138799;
		16'd1054 : result2 = 138846;
		16'd1055 : result2 = 138919;
		16'd1056 : result2 = 139018;
		16'd1057 : result2 = 139145;
		16'd1058 : result2 = 139300;
		16'd1059 : result2 = 139484;
		16'd1060 : result2 = 139697;
		16'd1061 : result2 = 139940;
		16'd1062 : result2 = 140214;
		16'd1063 : result2 = 140521;
		16'd1064 : result2 = 140860;
		16'd1065 : result2 = 141234;
		16'd1066 : result2 = 141644;
		16'd1067 : result2 = 142092;
		16'd1068 : result2 = 142578;
		16'd1069 : result2 = 143107;
		16'd1070 : result2 = 143679;
		16'd1071 : result2 = 144299;
		16'd1072 : result2 = 144970;
		16'd1073 : result2 = 145695;
		16'd1074 : result2 = 146482;
		16'd1280 : result2 = 141951;
		16'd1281 : result2 = 142021;
		16'd1282 : result2 = 142008;
		16'd1283 : result2 = 141926;
		16'd1284 : result2 = 141790;
		16'd1285 : result2 = 141610;
		16'd1286 : result2 = 141395;
		16'd1287 : result2 = 141155;
		16'd1288 : result2 = 140895;
		16'd1289 : result2 = 140623;
		16'd1290 : result2 = 140344;
		16'd1291 : result2 = 140061;
		16'd1292 : result2 = 139779;
		16'd1293 : result2 = 139502;
		16'd1294 : result2 = 139232;
		16'd1295 : result2 = 138972;
		16'd1296 : result2 = 138724;
		16'd1297 : result2 = 138489;
		16'd1298 : result2 = 138271;
		16'd1299 : result2 = 138069;
		16'd1300 : result2 = 137886;
		16'd1301 : result2 = 137723;
		16'd1302 : result2 = 137580;
		16'd1303 : result2 = 137458;
		16'd1304 : result2 = 137358;
		16'd1305 : result2 = 137281;
		16'd1306 : result2 = 137227;
		16'd1307 : result2 = 137198;
		16'd1308 : result2 = 137193;
		16'd1309 : result2 = 137213;
		16'd1310 : result2 = 137258;
		16'd1311 : result2 = 137330;
		16'd1312 : result2 = 137428;
		16'd1313 : result2 = 137553;
		16'd1314 : result2 = 137706;
		16'd1315 : result2 = 137887;
		16'd1316 : result2 = 138097;
		16'd1317 : result2 = 138337;
		16'd1318 : result2 = 138607;
		16'd1319 : result2 = 138909;
		16'd1320 : result2 = 139242;
		16'd1321 : result2 = 139610;
		16'd1322 : result2 = 140012;
		16'd1323 : result2 = 140451;
		16'd1324 : result2 = 140927;
		16'd1325 : result2 = 141444;
		16'd1326 : result2 = 142003;
		16'd1327 : result2 = 142607;
		16'd1328 : result2 = 143260;
		16'd1329 : result2 = 143965;
		16'd1330 : result2 = 144726;
		16'd1536 : result2 = 140133;
		16'd1537 : result2 = 140266;
		16'd1538 : result2 = 140300;
		16'd1539 : result2 = 140254;
		16'd1540 : result2 = 140144;
		16'd1541 : result2 = 139984;
		16'd1542 : result2 = 139785;
		16'd1543 : result2 = 139555;
		16'd1544 : result2 = 139304;
		16'd1545 : result2 = 139037;
		16'd1546 : result2 = 138761;
		16'd1547 : result2 = 138481;
		16'd1548 : result2 = 138201;
		16'd1549 : result2 = 137924;
		16'd1550 : result2 = 137655;
		16'd1551 : result2 = 137395;
		16'd1552 : result2 = 137146;
		16'd1553 : result2 = 136912;
		16'd1554 : result2 = 136693;
		16'd1555 : result2 = 136491;
		16'd1556 : result2 = 136308;
		16'd1557 : result2 = 136144;
		16'd1558 : result2 = 136001;
		16'd1559 : result2 = 135879;
		16'd1560 : result2 = 135779;
		16'd1561 : result2 = 135702;
		16'd1562 : result2 = 135648;
		16'd1563 : result2 = 135618;
		16'd1564 : result2 = 135613;
		16'd1565 : result2 = 135633;
		16'd1566 : result2 = 135678;
		16'd1567 : result2 = 135749;
		16'd1568 : result2 = 135846;
		16'd1569 : result2 = 135970;
		16'd1570 : result2 = 136122;
		16'd1571 : result2 = 136301;
		16'd1572 : result2 = 136509;
		16'd1573 : result2 = 136746;
		16'd1574 : result2 = 137014;
		16'd1575 : result2 = 137311;
		16'd1576 : result2 = 137641;
		16'd1577 : result2 = 138003;
		16'd1578 : result2 = 138399;
		16'd1579 : result2 = 138830;
		16'd1580 : result2 = 139298;
		16'd1581 : result2 = 139805;
		16'd1582 : result2 = 140353;
		16'd1583 : result2 = 140943;
		16'd1584 : result2 = 141580;
		16'd1585 : result2 = 142267;
		16'd1586 : result2 = 143007;
		16'd1792 : result2 = 138316;
		16'd1793 : result2 = 138516;
		16'd1794 : result2 = 138599;
		16'd1795 : result2 = 138590;
		16'd1796 : result2 = 138507;
		16'd1797 : result2 = 138367;
		16'd1798 : result2 = 138181;
		16'd1799 : result2 = 137962;
		16'd1800 : result2 = 137717;
		16'd1801 : result2 = 137456;
		16'd1802 : result2 = 137183;
		16'd1803 : result2 = 136905;
		16'd1804 : result2 = 136625;
		16'd1805 : result2 = 136349;
		16'd1806 : result2 = 136080;
		16'd1807 : result2 = 135820;
		16'd1808 : result2 = 135571;
		16'd1809 : result2 = 135336;
		16'd1810 : result2 = 135117;
		16'd1811 : result2 = 134915;
		16'd1812 : result2 = 134732;
		16'd1813 : result2 = 134568;
		16'd1814 : result2 = 134425;
		16'd1815 : result2 = 134303;
		16'd1816 : result2 = 134204;
		16'd1817 : result2 = 134127;
		16'd1818 : result2 = 134074;
		16'd1819 : result2 = 134044;
		16'd1820 : result2 = 134039;
		16'd1821 : result2 = 134059;
		16'd1822 : result2 = 134105;
		16'd1823 : result2 = 134176;
		16'd1824 : result2 = 134273;
		16'd1825 : result2 = 134397;
		16'd1826 : result2 = 134548;
		16'd1827 : result2 = 134726;
		16'd1828 : result2 = 134933;
		16'd1829 : result2 = 135168;
		16'd1830 : result2 = 135433;
		16'd1831 : result2 = 135728;
		16'd1832 : result2 = 136054;
		16'd1833 : result2 = 136412;
		16'd1834 : result2 = 136803;
		16'd1835 : result2 = 137228;
		16'd1836 : result2 = 137689;
		16'd1837 : result2 = 138187;
		16'd1838 : result2 = 138725;
		16'd1839 : result2 = 139305;
		16'd1840 : result2 = 139928;
		16'd1841 : result2 = 140599;
		16'd1842 : result2 = 141321;
		16'd2048 : result2 = 136506;
		16'd2049 : result2 = 136775;
		16'd2050 : result2 = 136909;
		16'd2051 : result2 = 136936;
		16'd2052 : result2 = 136880;
		16'd2053 : result2 = 136758;
		16'd2054 : result2 = 136586;
		16'd2055 : result2 = 136375;
		16'd2056 : result2 = 136137;
		16'd2057 : result2 = 135879;
		16'd2058 : result2 = 135608;
		16'd2059 : result2 = 135331;
		16'd2060 : result2 = 135053;
		16'd2061 : result2 = 134777;
		16'd2062 : result2 = 134507;
		16'd2063 : result2 = 134247;
		16'd2064 : result2 = 133998;
		16'd2065 : result2 = 133763;
		16'd2066 : result2 = 133543;
		16'd2067 : result2 = 133342;
		16'd2068 : result2 = 133158;
		16'd2069 : result2 = 132995;
		16'd2070 : result2 = 132852;
		16'd2071 : result2 = 132731;
		16'd2072 : result2 = 132632;
		16'd2073 : result2 = 132556;
		16'd2074 : result2 = 132503;
		16'd2075 : result2 = 132475;
		16'd2076 : result2 = 132471;
		16'd2077 : result2 = 132491;
		16'd2078 : result2 = 132537;
		16'd2079 : result2 = 132609;
		16'd2080 : result2 = 132707;
		16'd2081 : result2 = 132831;
		16'd2082 : result2 = 132982;
		16'd2083 : result2 = 133160;
		16'd2084 : result2 = 133366;
		16'd2085 : result2 = 133601;
		16'd2086 : result2 = 133864;
		16'd2087 : result2 = 134157;
		16'd2088 : result2 = 134481;
		16'd2089 : result2 = 134836;
		16'd2090 : result2 = 135223;
		16'd2091 : result2 = 135643;
		16'd2092 : result2 = 136098;
		16'd2093 : result2 = 136590;
		16'd2094 : result2 = 137119;
		16'd2095 : result2 = 137689;
		16'd2096 : result2 = 138301;
		16'd2097 : result2 = 138958;
		16'd2098 : result2 = 139664;
		16'd2304 : result2 = 134707;
		16'd2305 : result2 = 135049;
		16'd2306 : result2 = 135234;
		16'd2307 : result2 = 135297;
		16'd2308 : result2 = 135265;
		16'd2309 : result2 = 135160;
		16'd2310 : result2 = 134999;
		16'd2311 : result2 = 134796;
		16'd2312 : result2 = 134563;
		16'd2313 : result2 = 134307;
		16'd2314 : result2 = 134038;
		16'd2315 : result2 = 133762;
		16'd2316 : result2 = 133483;
		16'd2317 : result2 = 133207;
		16'd2318 : result2 = 132936;
		16'd2319 : result2 = 132675;
		16'd2320 : result2 = 132426;
		16'd2321 : result2 = 132190;
		16'd2322 : result2 = 131971;
		16'd2323 : result2 = 131769;
		16'd2324 : result2 = 131586;
		16'd2325 : result2 = 131423;
		16'd2326 : result2 = 131281;
		16'd2327 : result2 = 131160;
		16'd2328 : result2 = 131062;
		16'd2329 : result2 = 130988;
		16'd2330 : result2 = 130936;
		16'd2331 : result2 = 130909;
		16'd2332 : result2 = 130906;
		16'd2333 : result2 = 130928;
		16'd2334 : result2 = 130976;
		16'd2335 : result2 = 131049;
		16'd2336 : result2 = 131147;
		16'd2337 : result2 = 131273;
		16'd2338 : result2 = 131424;
		16'd2339 : result2 = 131603;
		16'd2340 : result2 = 131809;
		16'd2341 : result2 = 132044;
		16'd2342 : result2 = 132307;
		16'd2343 : result2 = 132599;
		16'd2344 : result2 = 132920;
		16'd2345 : result2 = 133273;
		16'd2346 : result2 = 133657;
		16'd2347 : result2 = 134074;
		16'd2348 : result2 = 134524;
		16'd2349 : result2 = 135010;
		16'd2350 : result2 = 135533;
		16'd2351 : result2 = 136094;
		16'd2352 : result2 = 136697;
		16'd2353 : result2 = 137343;
		16'd2354 : result2 = 138035;
		16'd2560 : result2 = 132928;
		16'd2561 : result2 = 133344;
		16'd2562 : result2 = 133578;
		16'd2563 : result2 = 133674;
		16'd2564 : result2 = 133665;
		16'd2565 : result2 = 133575;
		16'd2566 : result2 = 133424;
		16'd2567 : result2 = 133226;
		16'd2568 : result2 = 132996;
		16'd2569 : result2 = 132742;
		16'd2570 : result2 = 132473;
		16'd2571 : result2 = 132195;
		16'd2572 : result2 = 131916;
		16'd2573 : result2 = 131638;
		16'd2574 : result2 = 131367;
		16'd2575 : result2 = 131105;
		16'd2576 : result2 = 130854;
		16'd2577 : result2 = 130619;
		16'd2578 : result2 = 130399;
		16'd2579 : result2 = 130197;
		16'd2580 : result2 = 130015;
		16'd2581 : result2 = 129852;
		16'd2582 : result2 = 129711;
		16'd2583 : result2 = 129592;
		16'd2584 : result2 = 129495;
		16'd2585 : result2 = 129422;
		16'd2586 : result2 = 129372;
		16'd2587 : result2 = 129347;
		16'd2588 : result2 = 129346;
		16'd2589 : result2 = 129370;
		16'd2590 : result2 = 129419;
		16'd2591 : result2 = 129494;
		16'd2592 : result2 = 129594;
		16'd2593 : result2 = 129721;
		16'd2594 : result2 = 129874;
		16'd2595 : result2 = 130054;
		16'd2596 : result2 = 130261;
		16'd2597 : result2 = 130496;
		16'd2598 : result2 = 130759;
		16'd2599 : result2 = 131051;
		16'd2600 : result2 = 131372;
		16'd2601 : result2 = 131723;
		16'd2602 : result2 = 132105;
		16'd2603 : result2 = 132519;
		16'd2604 : result2 = 132967;
		16'd2605 : result2 = 133448;
		16'd2606 : result2 = 133965;
		16'd2607 : result2 = 134520;
		16'd2608 : result2 = 135114;
		16'd2609 : result2 = 135750;
		16'd2610 : result2 = 136431;
		16'd2816 : result2 = 131175;
		16'd2817 : result2 = 131664;
		16'd2818 : result2 = 131946;
		16'd2819 : result2 = 132073;
		16'd2820 : result2 = 132083;
		16'd2821 : result2 = 132005;
		16'd2822 : result2 = 131860;
		16'd2823 : result2 = 131666;
		16'd2824 : result2 = 131436;
		16'd2825 : result2 = 131182;
		16'd2826 : result2 = 130911;
		16'd2827 : result2 = 130632;
		16'd2828 : result2 = 130351;
		16'd2829 : result2 = 130072;
		16'd2830 : result2 = 129798;
		16'd2831 : result2 = 129535;
		16'd2832 : result2 = 129284;
		16'd2833 : result2 = 129047;
		16'd2834 : result2 = 128828;
		16'd2835 : result2 = 128626;
		16'd2836 : result2 = 128444;
		16'd2837 : result2 = 128282;
		16'd2838 : result2 = 128142;
		16'd2839 : result2 = 128025;
		16'd2840 : result2 = 127930;
		16'd2841 : result2 = 127858;
		16'd2842 : result2 = 127811;
		16'd2843 : result2 = 127788;
		16'd2844 : result2 = 127789;
		16'd2845 : result2 = 127815;
		16'd2846 : result2 = 127867;
		16'd2847 : result2 = 127944;
		16'd2848 : result2 = 128047;
		16'd2849 : result2 = 128175;
		16'd2850 : result2 = 128331;
		16'd2851 : result2 = 128512;
		16'd2852 : result2 = 128721;
		16'd2853 : result2 = 128957;
		16'd2854 : result2 = 129221;
		16'd2855 : result2 = 129513;
		16'd2856 : result2 = 129835;
		16'd2857 : result2 = 130185;
		16'd2858 : result2 = 130566;
		16'd2859 : result2 = 130979;
		16'd2860 : result2 = 131423;
		16'd2861 : result2 = 131901;
		16'd2862 : result2 = 132414;
		16'd2863 : result2 = 132964;
		16'd2864 : result2 = 133551;
		16'd2865 : result2 = 134179;
		16'd2866 : result2 = 134850;
		16'd3072 : result2 = 129459;
		16'd3073 : result2 = 130018;
		16'd3074 : result2 = 130342;
		16'd3075 : result2 = 130495;
		16'd3076 : result2 = 130521;
		16'd3077 : result2 = 130450;
		16'd3078 : result2 = 130309;
		16'd3079 : result2 = 130116;
		16'd3080 : result2 = 129884;
		16'd3081 : result2 = 129628;
		16'd3082 : result2 = 129355;
		16'd3083 : result2 = 129073;
		16'd3084 : result2 = 128788;
		16'd3085 : result2 = 128506;
		16'd3086 : result2 = 128231;
		16'd3087 : result2 = 127966;
		16'd3088 : result2 = 127713;
		16'd3089 : result2 = 127476;
		16'd3090 : result2 = 127256;
		16'd3091 : result2 = 127055;
		16'd3092 : result2 = 126873;
		16'd3093 : result2 = 126713;
		16'd3094 : result2 = 126574;
		16'd3095 : result2 = 126458;
		16'd3096 : result2 = 126365;
		16'd3097 : result2 = 126296;
		16'd3098 : result2 = 126251;
		16'd3099 : result2 = 126231;
		16'd3100 : result2 = 126235;
		16'd3101 : result2 = 126264;
		16'd3102 : result2 = 126319;
		16'd3103 : result2 = 126398;
		16'd3104 : result2 = 126504;
		16'd3105 : result2 = 126636;
		16'd3106 : result2 = 126793;
		16'd3107 : result2 = 126978;
		16'd3108 : result2 = 127188;
		16'd3109 : result2 = 127427;
		16'd3110 : result2 = 127692;
		16'd3111 : result2 = 127986;
		16'd3112 : result2 = 128308;
		16'd3113 : result2 = 128659;
		16'd3114 : result2 = 129040;
		16'd3115 : result2 = 129451;
		16'd3116 : result2 = 129894;
		16'd3117 : result2 = 130370;
		16'd3118 : result2 = 130879;
		16'd3119 : result2 = 131424;
		16'd3120 : result2 = 132006;
		16'd3121 : result2 = 132628;
		16'd3122 : result2 = 133290;
		16'd3328 : result2 = 127788;
		16'd3329 : result2 = 128411;
		16'd3330 : result2 = 128772;
		16'd3331 : result2 = 128945;
		16'd3332 : result2 = 128981;
		16'd3333 : result2 = 128914;
		16'd3334 : result2 = 128772;
		16'd3335 : result2 = 128576;
		16'd3336 : result2 = 128341;
		16'd3337 : result2 = 128080;
		16'd3338 : result2 = 127802;
		16'd3339 : result2 = 127516;
		16'd3340 : result2 = 127227;
		16'd3341 : result2 = 126942;
		16'd3342 : result2 = 126664;
		16'd3343 : result2 = 126397;
		16'd3344 : result2 = 126143;
		16'd3345 : result2 = 125905;
		16'd3346 : result2 = 125684;
		16'd3347 : result2 = 125483;
		16'd3348 : result2 = 125302;
		16'd3349 : result2 = 125143;
		16'd3350 : result2 = 125006;
		16'd3351 : result2 = 124892;
		16'd3352 : result2 = 124802;
		16'd3353 : result2 = 124735;
		16'd3354 : result2 = 124693;
		16'd3355 : result2 = 124676;
		16'd3356 : result2 = 124683;
		16'd3357 : result2 = 124716;
		16'd3358 : result2 = 124774;
		16'd3359 : result2 = 124857;
		16'd3360 : result2 = 124966;
		16'd3361 : result2 = 125101;
		16'd3362 : result2 = 125262;
		16'd3363 : result2 = 125449;
		16'd3364 : result2 = 125663;
		16'd3365 : result2 = 125903;
		16'd3366 : result2 = 126171;
		16'd3367 : result2 = 126467;
		16'd3368 : result2 = 126790;
		16'd3369 : result2 = 127142;
		16'd3370 : result2 = 127524;
		16'd3371 : result2 = 127935;
		16'd3372 : result2 = 128378;
		16'd3373 : result2 = 128852;
		16'd3374 : result2 = 129359;
		16'd3375 : result2 = 129901;
		16'd3376 : result2 = 130479;
		16'd3377 : result2 = 131095;
		16'd3378 : result2 = 131751;
		16'd3584 : result2 = 126173;
		16'd3585 : result2 = 126851;
		16'd3586 : result2 = 127241;
		16'd3587 : result2 = 127426;
		16'd3588 : result2 = 127465;
		16'd3589 : result2 = 127396;
		16'd3590 : result2 = 127250;
		16'd3591 : result2 = 127048;
		16'd3592 : result2 = 126806;
		16'd3593 : result2 = 126538;
		16'd3594 : result2 = 126253;
		16'd3595 : result2 = 125961;
		16'd3596 : result2 = 125668;
		16'd3597 : result2 = 125378;
		16'd3598 : result2 = 125097;
		16'd3599 : result2 = 124827;
		16'd3600 : result2 = 124571;
		16'd3601 : result2 = 124332;
		16'd3602 : result2 = 124111;
		16'd3603 : result2 = 123910;
		16'd3604 : result2 = 123731;
		16'd3605 : result2 = 123573;
		16'd3606 : result2 = 123438;
		16'd3607 : result2 = 123326;
		16'd3608 : result2 = 123239;
		16'd3609 : result2 = 123175;
		16'd3610 : result2 = 123137;
		16'd3611 : result2 = 123123;
		16'd3612 : result2 = 123134;
		16'd3613 : result2 = 123170;
		16'd3614 : result2 = 123232;
		16'd3615 : result2 = 123319;
		16'd3616 : result2 = 123432;
		16'd3617 : result2 = 123571;
		16'd3618 : result2 = 123736;
		16'd3619 : result2 = 123926;
		16'd3620 : result2 = 124144;
		16'd3621 : result2 = 124388;
		16'd3622 : result2 = 124658;
		16'd3623 : result2 = 124956;
		16'd3624 : result2 = 125282;
		16'd3625 : result2 = 125636;
		16'd3626 : result2 = 126019;
		16'd3627 : result2 = 126431;
		16'd3628 : result2 = 126874;
		16'd3629 : result2 = 127348;
		16'd3630 : result2 = 127854;
		16'd3631 : result2 = 128393;
		16'd3632 : result2 = 128968;
		16'd3633 : result2 = 129580;
		16'd3634 : result2 = 130230;
		16'd3840 : result2 = 124624;
		16'd3841 : result2 = 125345;
		16'd3842 : result2 = 125751;
		16'd3843 : result2 = 125940;
		16'd3844 : result2 = 125975;
		16'd3845 : result2 = 125899;
		16'd3846 : result2 = 125743;
		16'd3847 : result2 = 125530;
		16'd3848 : result2 = 125278;
		16'd3849 : result2 = 125001;
		16'd3850 : result2 = 124708;
		16'd3851 : result2 = 124409;
		16'd3852 : result2 = 124109;
		16'd3853 : result2 = 123814;
		16'd3854 : result2 = 123529;
		16'd3855 : result2 = 123256;
		16'd3856 : result2 = 122998;
		16'd3857 : result2 = 122758;
		16'd3858 : result2 = 122537;
		16'd3859 : result2 = 122336;
		16'd3860 : result2 = 122158;
		16'd3861 : result2 = 122002;
		16'd3862 : result2 = 121869;
		16'd3863 : result2 = 121760;
		16'd3864 : result2 = 121676;
		16'd3865 : result2 = 121616;
		16'd3866 : result2 = 121581;
		16'd3867 : result2 = 121571;
		16'd3868 : result2 = 121586;
		16'd3869 : result2 = 121627;
		16'd3870 : result2 = 121693;
		16'd3871 : result2 = 121785;
		16'd3872 : result2 = 121902;
		16'd3873 : result2 = 122045;
		16'd3874 : result2 = 122214;
		16'd3875 : result2 = 122409;
		16'd3876 : result2 = 122631;
		16'd3877 : result2 = 122878;
		16'd3878 : result2 = 123153;
		16'd3879 : result2 = 123454;
		16'd3880 : result2 = 123783;
		16'd3881 : result2 = 124139;
		16'd3882 : result2 = 124524;
		16'd3883 : result2 = 124938;
		16'd3884 : result2 = 125381;
		16'd3885 : result2 = 125855;
		16'd3886 : result2 = 126361;
		16'd3887 : result2 = 126900;
		16'd3888 : result2 = 127472;
		16'd3889 : result2 = 128081;
		16'd3890 : result2 = 128727;
		16'd4096 : result2 = 123151;
		16'd4097 : result2 = 123897;
		16'd4098 : result2 = 124307;
		16'd4099 : result2 = 124488;
		16'd4100 : result2 = 124511;
		16'd4101 : result2 = 124420;
		16'd4102 : result2 = 124250;
		16'd4103 : result2 = 124023;
		16'd4104 : result2 = 123758;
		16'd4105 : result2 = 123469;
		16'd4106 : result2 = 123166;
		16'd4107 : result2 = 122857;
		16'd4108 : result2 = 122550;
		16'd4109 : result2 = 122250;
		16'd4110 : result2 = 121959;
		16'd4111 : result2 = 121683;
		16'd4112 : result2 = 121423;
		16'd4113 : result2 = 121181;
		16'd4114 : result2 = 120960;
		16'd4115 : result2 = 120760;
		16'd4116 : result2 = 120583;
		16'd4117 : result2 = 120429;
		16'd4118 : result2 = 120299;
		16'd4119 : result2 = 120193;
		16'd4120 : result2 = 120112;
		16'd4121 : result2 = 120056;
		16'd4122 : result2 = 120025;
		16'd4123 : result2 = 120020;
		16'd4124 : result2 = 120040;
		16'd4125 : result2 = 120086;
		16'd4126 : result2 = 120157;
		16'd4127 : result2 = 120253;
		16'd4128 : result2 = 120376;
		16'd4129 : result2 = 120524;
		16'd4130 : result2 = 120698;
		16'd4131 : result2 = 120898;
		16'd4132 : result2 = 121123;
		16'd4133 : result2 = 121375;
		16'd4134 : result2 = 121654;
		16'd4135 : result2 = 121959;
		16'd4136 : result2 = 122291;
		16'd4137 : result2 = 122651;
		16'd4138 : result2 = 123039;
		16'd4139 : result2 = 123455;
		16'd4140 : result2 = 123900;
		16'd4141 : result2 = 124375;
		16'd4142 : result2 = 124881;
		16'd4143 : result2 = 125420;
		16'd4144 : result2 = 125991;
		16'd4145 : result2 = 126597;
		16'd4146 : result2 = 127240;
		16'd4352 : result2 = 121763;
		16'd4353 : result2 = 122512;
		16'd4354 : result2 = 122909;
		16'd4355 : result2 = 123072;
		16'd4356 : result2 = 123073;
		16'd4357 : result2 = 122961;
		16'd4358 : result2 = 122770;
		16'd4359 : result2 = 122525;
		16'd4360 : result2 = 122244;
		16'd4361 : result2 = 121940;
		16'd4362 : result2 = 121625;
		16'd4363 : result2 = 121307;
		16'd4364 : result2 = 120991;
		16'd4365 : result2 = 120683;
		16'd4366 : result2 = 120388;
		16'd4367 : result2 = 120108;
		16'd4368 : result2 = 119845;
		16'd4369 : result2 = 119602;
		16'd4370 : result2 = 119381;
		16'd4371 : result2 = 119182;
		16'd4372 : result2 = 119006;
		16'd4373 : result2 = 118854;
		16'd4374 : result2 = 118727;
		16'd4375 : result2 = 118625;
		16'd4376 : result2 = 118548;
		16'd4377 : result2 = 118496;
		16'd4378 : result2 = 118470;
		16'd4379 : result2 = 118470;
		16'd4380 : result2 = 118495;
		16'd4381 : result2 = 118546;
		16'd4382 : result2 = 118622;
		16'd4383 : result2 = 118725;
		16'd4384 : result2 = 118852;
		16'd4385 : result2 = 119006;
		16'd4386 : result2 = 119185;
		16'd4387 : result2 = 119391;
		16'd4388 : result2 = 119622;
		16'd4389 : result2 = 119879;
		16'd4390 : result2 = 120162;
		16'd4391 : result2 = 120472;
		16'd4392 : result2 = 120808;
		16'd4393 : result2 = 121171;
		16'd4394 : result2 = 121562;
		16'd4395 : result2 = 121981;
		16'd4396 : result2 = 122429;
		16'd4397 : result2 = 122906;
		16'd4398 : result2 = 123414;
		16'd4399 : result2 = 123952;
		16'd4400 : result2 = 124524;
		16'd4401 : result2 = 125129;
		16'd4402 : result2 = 125769;
		16'd4608 : result2 = 120464;
		16'd4609 : result2 = 121193;
		16'd4610 : result2 = 121560;
		16'd4611 : result2 = 121691;
		16'd4612 : result2 = 121661;
		16'd4613 : result2 = 121520;
		16'd4614 : result2 = 121304;
		16'd4615 : result2 = 121036;
		16'd4616 : result2 = 120735;
		16'd4617 : result2 = 120415;
		16'd4618 : result2 = 120085;
		16'd4619 : result2 = 119755;
		16'd4620 : result2 = 119430;
		16'd4621 : result2 = 119115;
		16'd4622 : result2 = 118814;
		16'd4623 : result2 = 118529;
		16'd4624 : result2 = 118264;
		16'd4625 : result2 = 118020;
		16'd4626 : result2 = 117799;
		16'd4627 : result2 = 117600;
		16'd4628 : result2 = 117426;
		16'd4629 : result2 = 117277;
		16'd4630 : result2 = 117153;
		16'd4631 : result2 = 117055;
		16'd4632 : result2 = 116982;
		16'd4633 : result2 = 116935;
		16'd4634 : result2 = 116914;
		16'd4635 : result2 = 116919;
		16'd4636 : result2 = 116950;
		16'd4637 : result2 = 117007;
		16'd4638 : result2 = 117090;
		16'd4639 : result2 = 117198;
		16'd4640 : result2 = 117332;
		16'd4641 : result2 = 117492;
		16'd4642 : result2 = 117677;
		16'd4643 : result2 = 117888;
		16'd4644 : result2 = 118125;
		16'd4645 : result2 = 118388;
		16'd4646 : result2 = 118676;
		16'd4647 : result2 = 118991;
		16'd4648 : result2 = 119332;
		16'd4649 : result2 = 119700;
		16'd4650 : result2 = 120095;
		16'd4651 : result2 = 120517;
		16'd4652 : result2 = 120968;
		16'd4653 : result2 = 121448;
		16'd4654 : result2 = 121957;
		16'd4655 : result2 = 122497;
		16'd4656 : result2 = 123069;
		16'd4657 : result2 = 123674;
		16'd4658 : result2 = 124314;
		16'd4864 : result2 = 119257;
		16'd4865 : result2 = 119938;
		16'd4866 : result2 = 120256;
		16'd4867 : result2 = 120342;
		16'd4868 : result2 = 120271;
		16'd4869 : result2 = 120095;
		16'd4870 : result2 = 119847;
		16'd4871 : result2 = 119553;
		16'd4872 : result2 = 119229;
		16'd4873 : result2 = 118890;
		16'd4874 : result2 = 118545;
		16'd4875 : result2 = 118201;
		16'd4876 : result2 = 117866;
		16'd4877 : result2 = 117543;
		16'd4878 : result2 = 117236;
		16'd4879 : result2 = 116947;
		16'd4880 : result2 = 116679;
		16'd4881 : result2 = 116434;
		16'd4882 : result2 = 116212;
		16'd4883 : result2 = 116015;
		16'd4884 : result2 = 115843;
		16'd4885 : result2 = 115697;
		16'd4886 : result2 = 115577;
		16'd4887 : result2 = 115483;
		16'd4888 : result2 = 115415;
		16'd4889 : result2 = 115374;
		16'd4890 : result2 = 115358;
		16'd4891 : result2 = 115370;
		16'd4892 : result2 = 115407;
		16'd4893 : result2 = 115470;
		16'd4894 : result2 = 115559;
		16'd4895 : result2 = 115674;
		16'd4896 : result2 = 115815;
		16'd4897 : result2 = 115981;
		16'd4898 : result2 = 116173;
		16'd4899 : result2 = 116390;
		16'd4900 : result2 = 116633;
		16'd4901 : result2 = 116902;
		16'd4902 : result2 = 117196;
		16'd4903 : result2 = 117517;
		16'd4904 : result2 = 117863;
		16'd4905 : result2 = 118236;
		16'd4906 : result2 = 118636;
		16'd4907 : result2 = 119063;
		16'd4908 : result2 = 119517;
		16'd4909 : result2 = 120000;
		16'd4910 : result2 = 120512;
		16'd4911 : result2 = 121054;
		16'd4912 : result2 = 121627;
		16'd4913 : result2 = 122233;
		16'd4914 : result2 = 122872;
		16'd5120 : result2 = 118140;
		16'd5121 : result2 = 118744;
		16'd5122 : result2 = 118995;
		16'd5123 : result2 = 119022;
		16'd5124 : result2 = 118902;
		16'd5125 : result2 = 118683;
		16'd5126 : result2 = 118399;
		16'd5127 : result2 = 118074;
		16'd5128 : result2 = 117725;
		16'd5129 : result2 = 117364;
		16'd5130 : result2 = 117002;
		16'd5131 : result2 = 116644;
		16'd5132 : result2 = 116298;
		16'd5133 : result2 = 115966;
		16'd5134 : result2 = 115653;
		16'd5135 : result2 = 115360;
		16'd5136 : result2 = 115090;
		16'd5137 : result2 = 114843;
		16'd5138 : result2 = 114622;
		16'd5139 : result2 = 114426;
		16'd5140 : result2 = 114257;
		16'd5141 : result2 = 114114;
		16'd5142 : result2 = 113998;
		16'd5143 : result2 = 113909;
		16'd5144 : result2 = 113846;
		16'd5145 : result2 = 113811;
		16'd5146 : result2 = 113802;
		16'd5147 : result2 = 113819;
		16'd5148 : result2 = 113863;
		16'd5149 : result2 = 113933;
		16'd5150 : result2 = 114030;
		16'd5151 : result2 = 114152;
		16'd5152 : result2 = 114300;
		16'd5153 : result2 = 114473;
		16'd5154 : result2 = 114672;
		16'd5155 : result2 = 114896;
		16'd5156 : result2 = 115146;
		16'd5157 : result2 = 115422;
		16'd5158 : result2 = 115723;
		16'd5159 : result2 = 116049;
		16'd5160 : result2 = 116402;
		16'd5161 : result2 = 116780;
		16'd5162 : result2 = 117185;
		16'd5163 : result2 = 117617;
		16'd5164 : result2 = 118075;
		16'd5165 : result2 = 118562;
		16'd5166 : result2 = 119078;
		16'd5167 : result2 = 119622;
		16'd5168 : result2 = 120198;
		16'd5169 : result2 = 120804;
		16'd5170 : result2 = 121444;
		16'd5376 : result2 = 117105;
		16'd5377 : result2 = 117605;
		16'd5378 : result2 = 117770;
		16'd5379 : result2 = 117727;
		16'd5380 : result2 = 117547;
		16'd5381 : result2 = 117280;
		16'd5382 : result2 = 116955;
		16'd5383 : result2 = 116597;
		16'd5384 : result2 = 116220;
		16'd5385 : result2 = 115836;
		16'd5386 : result2 = 115455;
		16'd5387 : result2 = 115083;
		16'd5388 : result2 = 114724;
		16'd5389 : result2 = 114384;
		16'd5390 : result2 = 114064;
		16'd5391 : result2 = 113767;
		16'd5392 : result2 = 113494;
		16'd5393 : result2 = 113247;
		16'd5394 : result2 = 113027;
		16'd5395 : result2 = 112833;
		16'd5396 : result2 = 112666;
		16'd5397 : result2 = 112527;
		16'd5398 : result2 = 112416;
		16'd5399 : result2 = 112332;
		16'd5400 : result2 = 112276;
		16'd5401 : result2 = 112246;
		16'd5402 : result2 = 112244;
		16'd5403 : result2 = 112269;
		16'd5404 : result2 = 112320;
		16'd5405 : result2 = 112398;
		16'd5406 : result2 = 112502;
		16'd5407 : result2 = 112631;
		16'd5408 : result2 = 112787;
		16'd5409 : result2 = 112968;
		16'd5410 : result2 = 113175;
		16'd5411 : result2 = 113407;
		16'd5412 : result2 = 113664;
		16'd5413 : result2 = 113947;
		16'd5414 : result2 = 114254;
		16'd5415 : result2 = 114588;
		16'd5416 : result2 = 114947;
		16'd5417 : result2 = 115331;
		16'd5418 : result2 = 115742;
		16'd5419 : result2 = 116179;
		16'd5420 : result2 = 116643;
		16'd5421 : result2 = 117134;
		16'd5422 : result2 = 117654;
		16'd5423 : result2 = 118202;
		16'd5424 : result2 = 118780;
		16'd5425 : result2 = 119389;
		16'd5426 : result2 = 120030;
		16'd5632 : result2 = 116141;
		16'd5633 : result2 = 116510;
		16'd5634 : result2 = 116574;
		16'd5635 : result2 = 116449;
		16'd5636 : result2 = 116204;
		16'd5637 : result2 = 115882;
		16'd5638 : result2 = 115513;
		16'd5639 : result2 = 115117;
		16'd5640 : result2 = 114710;
		16'd5641 : result2 = 114303;
		16'd5642 : result2 = 113902;
		16'd5643 : result2 = 113514;
		16'd5644 : result2 = 113144;
		16'd5645 : result2 = 112794;
		16'd5646 : result2 = 112468;
		16'd5647 : result2 = 112167;
		16'd5648 : result2 = 111892;
		16'd5649 : result2 = 111645;
		16'd5650 : result2 = 111425;
		16'd5651 : result2 = 111234;
		16'd5652 : result2 = 111071;
		16'd5653 : result2 = 110937;
		16'd5654 : result2 = 110830;
		16'd5655 : result2 = 110752;
		16'd5656 : result2 = 110702;
		16'd5657 : result2 = 110680;
		16'd5658 : result2 = 110685;
		16'd5659 : result2 = 110718;
		16'd5660 : result2 = 110777;
		16'd5661 : result2 = 110863;
		16'd5662 : result2 = 110975;
		16'd5663 : result2 = 111113;
		16'd5664 : result2 = 111277;
		16'd5665 : result2 = 111466;
		16'd5666 : result2 = 111681;
		16'd5667 : result2 = 111921;
		16'd5668 : result2 = 112186;
		16'd5669 : result2 = 112476;
		16'd5670 : result2 = 112792;
		16'd5671 : result2 = 113132;
		16'd5672 : result2 = 113498;
		16'd5673 : result2 = 113890;
		16'd5674 : result2 = 114307;
		16'd5675 : result2 = 114750;
		16'd5676 : result2 = 115219;
		16'd5677 : result2 = 115716;
		16'd5678 : result2 = 116239;
		16'd5679 : result2 = 116792;
		16'd5680 : result2 = 117373;
		16'd5681 : result2 = 117985;
		16'd5682 : result2 = 118628;
		16'd5888 : result2 = 115229;
		16'd5889 : result2 = 115448;
		16'd5890 : result2 = 115397;
		16'd5891 : result2 = 115182;
		16'd5892 : result2 = 114864;
		16'd5893 : result2 = 114484;
		16'd5894 : result2 = 114067;
		16'd5895 : result2 = 113633;
		16'd5896 : result2 = 113195;
		16'd5897 : result2 = 112761;
		16'd5898 : result2 = 112341;
		16'd5899 : result2 = 111937;
		16'd5900 : result2 = 111555;
		16'd5901 : result2 = 111197;
		16'd5902 : result2 = 110865;
		16'd5903 : result2 = 110560;
		16'd5904 : result2 = 110283;
		16'd5905 : result2 = 110036;
		16'd5906 : result2 = 109818;
		16'd5907 : result2 = 109630;
		16'd5908 : result2 = 109471;
		16'd5909 : result2 = 109342;
		16'd5910 : result2 = 109241;
		16'd5911 : result2 = 109170;
		16'd5912 : result2 = 109127;
		16'd5913 : result2 = 109112;
		16'd5914 : result2 = 109125;
		16'd5915 : result2 = 109166;
		16'd5916 : result2 = 109234;
		16'd5917 : result2 = 109328;
		16'd5918 : result2 = 109449;
		16'd5919 : result2 = 109596;
		16'd5920 : result2 = 109768;
		16'd5921 : result2 = 109967;
		16'd5922 : result2 = 110190;
		16'd5923 : result2 = 110439;
		16'd5924 : result2 = 110713;
		16'd5925 : result2 = 111011;
		16'd5926 : result2 = 111335;
		16'd5927 : result2 = 111683;
		16'd5928 : result2 = 112057;
		16'd5929 : result2 = 112455;
		16'd5930 : result2 = 112879;
		16'd5931 : result2 = 113329;
		16'd5932 : result2 = 113804;
		16'd5933 : result2 = 114306;
		16'd5934 : result2 = 114835;
		16'd5935 : result2 = 115392;
		16'd5936 : result2 = 115978;
		16'd5937 : result2 = 116593;
		16'd5938 : result2 = 117238;
		16'd6144 : result2 = 114351;
		16'd6145 : result2 = 114404;
		16'd6146 : result2 = 114229;
		16'd6147 : result2 = 113917;
		16'd6148 : result2 = 113522;
		16'd6149 : result2 = 113080;
		16'd6150 : result2 = 112614;
		16'd6151 : result2 = 112140;
		16'd6152 : result2 = 111669;
		16'd6153 : result2 = 111210;
		16'd6154 : result2 = 110769;
		16'd6155 : result2 = 110350;
		16'd6156 : result2 = 109956;
		16'd6157 : result2 = 109589;
		16'd6158 : result2 = 109252;
		16'd6159 : result2 = 108944;
		16'd6160 : result2 = 108666;
		16'd6161 : result2 = 108420;
		16'd6162 : result2 = 108204;
		16'd6163 : result2 = 108019;
		16'd6164 : result2 = 107865;
		16'd6165 : result2 = 107742;
		16'd6166 : result2 = 107648;
		16'd6167 : result2 = 107584;
		16'd6168 : result2 = 107548;
		16'd6169 : result2 = 107542;
		16'd6170 : result2 = 107564;
		16'd6171 : result2 = 107613;
		16'd6172 : result2 = 107690;
		16'd6173 : result2 = 107794;
		16'd6174 : result2 = 107924;
		16'd6175 : result2 = 108080;
		16'd6176 : result2 = 108262;
		16'd6177 : result2 = 108470;
		16'd6178 : result2 = 108703;
		16'd6179 : result2 = 108961;
		16'd6180 : result2 = 109243;
		16'd6181 : result2 = 109551;
		16'd6182 : result2 = 109883;
		16'd6183 : result2 = 110240;
		16'd6184 : result2 = 110621;
		16'd6185 : result2 = 111028;
		16'd6186 : result2 = 111459;
		16'd6187 : result2 = 111915;
		16'd6188 : result2 = 112398;
		16'd6189 : result2 = 112906;
		16'd6190 : result2 = 113441;
		16'd6191 : result2 = 114003;
		16'd6192 : result2 = 114593;
		16'd6193 : result2 = 115212;
		16'd6194 : result2 = 115861;
		16'd6400 : result2 = 113485;
		16'd6401 : result2 = 113363;
		16'd6402 : result2 = 113057;
		16'd6403 : result2 = 112644;
		16'd6404 : result2 = 112170;
		16'd6405 : result2 = 111665;
		16'd6406 : result2 = 111148;
		16'd6407 : result2 = 110633;
		16'd6408 : result2 = 110130;
		16'd6409 : result2 = 109646;
		16'd6410 : result2 = 109185;
		16'd6411 : result2 = 108750;
		16'd6412 : result2 = 108345;
		16'd6413 : result2 = 107971;
		16'd6414 : result2 = 107628;
		16'd6415 : result2 = 107318;
		16'd6416 : result2 = 107040;
		16'd6417 : result2 = 106795;
		16'd6418 : result2 = 106583;
		16'd6419 : result2 = 106402;
		16'd6420 : result2 = 106254;
		16'd6421 : result2 = 106137;
		16'd6422 : result2 = 106050;
		16'd6423 : result2 = 105994;
		16'd6424 : result2 = 105967;
		16'd6425 : result2 = 105970;
		16'd6426 : result2 = 106001;
		16'd6427 : result2 = 106060;
		16'd6428 : result2 = 106146;
		16'd6429 : result2 = 106260;
		16'd6430 : result2 = 106400;
		16'd6431 : result2 = 106567;
		16'd6432 : result2 = 106759;
		16'd6433 : result2 = 106976;
		16'd6434 : result2 = 107219;
		16'd6435 : result2 = 107486;
		16'd6436 : result2 = 107779;
		16'd6437 : result2 = 108095;
		16'd6438 : result2 = 108437;
		16'd6439 : result2 = 108802;
		16'd6440 : result2 = 109192;
		16'd6441 : result2 = 109607;
		16'd6442 : result2 = 110046;
		16'd6443 : result2 = 110510;
		16'd6444 : result2 = 110999;
		16'd6445 : result2 = 111514;
		16'd6446 : result2 = 112055;
		16'd6447 : result2 = 112623;
		16'd6448 : result2 = 113219;
		16'd6449 : result2 = 113842;
		16'd6450 : result2 = 114496;
		16'd6656 : result2 = 112607;
		16'd6657 : result2 = 112307;
		16'd6658 : result2 = 111869;
		16'd6659 : result2 = 111354;
		16'd6660 : result2 = 110800;
		16'd6661 : result2 = 110232;
		16'd6662 : result2 = 109665;
		16'd6663 : result2 = 109110;
		16'd6664 : result2 = 108575;
		16'd6665 : result2 = 108066;
		16'd6666 : result2 = 107586;
		16'd6667 : result2 = 107137;
		16'd6668 : result2 = 106721;
		16'd6669 : result2 = 106340;
		16'd6670 : result2 = 105993;
		16'd6671 : result2 = 105682;
		16'd6672 : result2 = 105405;
		16'd6673 : result2 = 105162;
		16'd6674 : result2 = 104953;
		16'd6675 : result2 = 104778;
		16'd6676 : result2 = 104636;
		16'd6677 : result2 = 104526;
		16'd6678 : result2 = 104448;
		16'd6679 : result2 = 104400;
		16'd6680 : result2 = 104383;
		16'd6681 : result2 = 104395;
		16'd6682 : result2 = 104436;
		16'd6683 : result2 = 104505;
		16'd6684 : result2 = 104602;
		16'd6685 : result2 = 104726;
		16'd6686 : result2 = 104877;
		16'd6687 : result2 = 105054;
		16'd6688 : result2 = 105257;
		16'd6689 : result2 = 105485;
		16'd6690 : result2 = 105738;
		16'd6691 : result2 = 106016;
		16'd6692 : result2 = 106318;
		16'd6693 : result2 = 106645;
		16'd6694 : result2 = 106996;
		16'd6695 : result2 = 107371;
		16'd6696 : result2 = 107770;
		16'd6697 : result2 = 108193;
		16'd6698 : result2 = 108641;
		16'd6699 : result2 = 109113;
		16'd6700 : result2 = 109610;
		16'd6701 : result2 = 110132;
		16'd6702 : result2 = 110680;
		16'd6703 : result2 = 111254;
		16'd6704 : result2 = 111855;
		16'd6705 : result2 = 112484;
		16'd6706 : result2 = 113142;
		16'd6912 : result2 = 111696;
		16'd6913 : result2 = 111222;
		16'd6914 : result2 = 110654;
		16'd6915 : result2 = 110039;
		16'd6916 : result2 = 109406;
		16'd6917 : result2 = 108776;
		16'd6918 : result2 = 108159;
		16'd6919 : result2 = 107566;
		16'd6920 : result2 = 107000;
		16'd6921 : result2 = 106467;
		16'd6922 : result2 = 105969;
		16'd6923 : result2 = 105507;
		16'd6924 : result2 = 105082;
		16'd6925 : result2 = 104695;
		16'd6926 : result2 = 104346;
		16'd6927 : result2 = 104034;
		16'd6928 : result2 = 103758;
		16'd6929 : result2 = 103519;
		16'd6930 : result2 = 103316;
		16'd6931 : result2 = 103147;
		16'd6932 : result2 = 103012;
		16'd6933 : result2 = 102910;
		16'd6934 : result2 = 102840;
		16'd6935 : result2 = 102802;
		16'd6936 : result2 = 102795;
		16'd6937 : result2 = 102818;
		16'd6938 : result2 = 102870;
		16'd6939 : result2 = 102950;
		16'd6940 : result2 = 103058;
		16'd6941 : result2 = 103193;
		16'd6942 : result2 = 103355;
		16'd6943 : result2 = 103544;
		16'd6944 : result2 = 103757;
		16'd6945 : result2 = 103997;
		16'd6946 : result2 = 104261;
		16'd6947 : result2 = 104549;
		16'd6948 : result2 = 104862;
		16'd6949 : result2 = 105199;
		16'd6950 : result2 = 105560;
		16'd6951 : result2 = 105945;
		16'd6952 : result2 = 106353;
		16'd6953 : result2 = 106786;
		16'd6954 : result2 = 107242;
		16'd6955 : result2 = 107723;
		16'd6956 : result2 = 108228;
		16'd6957 : result2 = 108758;
		16'd6958 : result2 = 109313;
		16'd6959 : result2 = 109894;
		16'd6960 : result2 = 110501;
		16'd6961 : result2 = 111136;
		16'd6962 : result2 = 111799;
		16'd7168 : result2 = 110733;
		16'd7169 : result2 = 110093;
		16'd7170 : result2 = 109400;
		16'd7171 : result2 = 108688;
		16'd7172 : result2 = 107981;
		16'd7173 : result2 = 107290;
		16'd7174 : result2 = 106627;
		16'd7175 : result2 = 105996;
		16'd7176 : result2 = 105402;
		16'd7177 : result2 = 104847;
		16'd7178 : result2 = 104333;
		16'd7179 : result2 = 103859;
		16'd7180 : result2 = 103427;
		16'd7181 : result2 = 103036;
		16'd7182 : result2 = 102684;
		16'd7183 : result2 = 102373;
		16'd7184 : result2 = 102101;
		16'd7185 : result2 = 101866;
		16'd7186 : result2 = 101669;
		16'd7187 : result2 = 101507;
		16'd7188 : result2 = 101381;
		16'd7189 : result2 = 101288;
		16'd7190 : result2 = 101228;
		16'd7191 : result2 = 101201;
		16'd7192 : result2 = 101204;
		16'd7193 : result2 = 101238;
		16'd7194 : result2 = 101301;
		16'd7195 : result2 = 101393;
		16'd7196 : result2 = 101513;
		16'd7197 : result2 = 101661;
		16'd7198 : result2 = 101835;
		16'd7199 : result2 = 102035;
		16'd7200 : result2 = 102260;
		16'd7201 : result2 = 102511;
		16'd7202 : result2 = 102786;
		16'd7203 : result2 = 103086;
		16'd7204 : result2 = 103410;
		16'd7205 : result2 = 103758;
		16'd7206 : result2 = 104130;
		16'd7207 : result2 = 104525;
		16'd7208 : result2 = 104944;
		16'd7209 : result2 = 105386;
		16'd7210 : result2 = 105852;
		16'd7211 : result2 = 106341;
		16'd7212 : result2 = 106855;
		16'd7213 : result2 = 107393;
		16'd7214 : result2 = 107956;
		16'd7215 : result2 = 108544;
		16'd7216 : result2 = 109158;
		16'd7217 : result2 = 109799;
		16'd7218 : result2 = 110468;
		16'd7424 : result2 = 109701;
		16'd7425 : result2 = 108907;
		16'd7426 : result2 = 108097;
		16'd7427 : result2 = 107295;
		16'd7428 : result2 = 106517;
		16'd7429 : result2 = 105771;
		16'd7430 : result2 = 105064;
		16'd7431 : result2 = 104399;
		16'd7432 : result2 = 103779;
		16'd7433 : result2 = 103204;
		16'd7434 : result2 = 102675;
		16'd7435 : result2 = 102192;
		16'd7436 : result2 = 101754;
		16'd7437 : result2 = 101359;
		16'd7438 : result2 = 101008;
		16'd7439 : result2 = 100699;
		16'd7440 : result2 = 100431;
		16'd7441 : result2 = 100203;
		16'd7442 : result2 = 100013;
		16'd7443 : result2 = 99859;
		16'd7444 : result2 = 99742;
		16'd7445 : result2 = 99660;
		16'd7446 : result2 = 99611;
		16'd7447 : result2 = 99595;
		16'd7448 : result2 = 99610;
		16'd7449 : result2 = 99656;
		16'd7450 : result2 = 99732;
		16'd7451 : result2 = 99836;
		16'd7452 : result2 = 99969;
		16'd7453 : result2 = 100128;
		16'd7454 : result2 = 100315;
		16'd7455 : result2 = 100527;
		16'd7456 : result2 = 100765;
		16'd7457 : result2 = 101028;
		16'd7458 : result2 = 101316;
		16'd7459 : result2 = 101628;
		16'd7460 : result2 = 101963;
		16'd7461 : result2 = 102323;
		16'd7462 : result2 = 102705;
		16'd7463 : result2 = 103111;
		16'd7464 : result2 = 103540;
		16'd7465 : result2 = 103993;
		16'd7466 : result2 = 104468;
		16'd7467 : result2 = 104967;
		16'd7468 : result2 = 105490;
		16'd7469 : result2 = 106037;
		16'd7470 : result2 = 106608;
		16'd7471 : result2 = 107204;
		16'd7472 : result2 = 107825;
		16'd7473 : result2 = 108473;
		16'd7474 : result2 = 109147;
		16'd7680 : result2 = 108586;
		16'd7681 : result2 = 107653;
		16'd7682 : result2 = 106736;
		16'd7683 : result2 = 105851;
		16'd7684 : result2 = 105008;
		16'd7685 : result2 = 104211;
		16'd7686 : result2 = 103465;
		16'd7687 : result2 = 102769;
		16'd7688 : result2 = 102126;
		16'd7689 : result2 = 101534;
		16'd7690 : result2 = 100994;
		16'd7691 : result2 = 100503;
		16'd7692 : result2 = 100061;
		16'd7693 : result2 = 99666;
		16'd7694 : result2 = 99317;
		16'd7695 : result2 = 99012;
		16'd7696 : result2 = 98749;
		16'd7697 : result2 = 98528;
		16'd7698 : result2 = 98347;
		16'd7699 : result2 = 98203;
		16'd7700 : result2 = 98097;
		16'd7701 : result2 = 98026;
		16'd7702 : result2 = 97989;
		16'd7703 : result2 = 97985;
		16'd7704 : result2 = 98013;
		16'd7705 : result2 = 98072;
		16'd7706 : result2 = 98160;
		16'd7707 : result2 = 98278;
		16'd7708 : result2 = 98424;
		16'd7709 : result2 = 98597;
		16'd7710 : result2 = 98796;
		16'd7711 : result2 = 99022;
		16'd7712 : result2 = 99273;
		16'd7713 : result2 = 99549;
		16'd7714 : result2 = 99849;
		16'd7715 : result2 = 100173;
		16'd7716 : result2 = 100521;
		16'd7717 : result2 = 100892;
		16'd7718 : result2 = 101286;
		16'd7719 : result2 = 101703;
		16'd7720 : result2 = 102143;
		16'd7721 : result2 = 102606;
		16'd7722 : result2 = 103092;
		16'd7723 : result2 = 103601;
		16'd7724 : result2 = 104133;
		16'd7725 : result2 = 104689;
		16'd7726 : result2 = 105269;
		16'd7727 : result2 = 105873;
		16'd7728 : result2 = 106502;
		16'd7729 : result2 = 107157;
		16'd7730 : result2 = 107838;
		16'd7936 : result2 = 107376;
		16'd7937 : result2 = 106321;
		16'd7938 : result2 = 105310;
		16'd7939 : result2 = 104351;
		16'd7940 : result2 = 103450;
		16'd7941 : result2 = 102608;
		16'd7942 : result2 = 101827;
		16'd7943 : result2 = 101105;
		16'd7944 : result2 = 100442;
		16'd7945 : result2 = 99837;
		16'd7946 : result2 = 99287;
		16'd7947 : result2 = 98791;
		16'd7948 : result2 = 98348;
		16'd7949 : result2 = 97954;
		16'd7950 : result2 = 97609;
		16'd7951 : result2 = 97310;
		16'd7952 : result2 = 97055;
		16'd7953 : result2 = 96842;
		16'd7954 : result2 = 96671;
		16'd7955 : result2 = 96538;
		16'd7956 : result2 = 96444;
		16'd7957 : result2 = 96385;
		16'd7958 : result2 = 96361;
		16'd7959 : result2 = 96371;
		16'd7960 : result2 = 96412;
		16'd7961 : result2 = 96485;
		16'd7962 : result2 = 96588;
		16'd7963 : result2 = 96719;
		16'd7964 : result2 = 96879;
		16'd7965 : result2 = 97066;
		16'd7966 : result2 = 97280;
		16'd7967 : result2 = 97519;
		16'd7968 : result2 = 97784;
		16'd7969 : result2 = 98073;
		16'd7970 : result2 = 98386;
		16'd7971 : result2 = 98723;
		16'd7972 : result2 = 99083;
		16'd7973 : result2 = 99467;
		16'd7974 : result2 = 99873;
		16'd7975 : result2 = 100302;
		16'd7976 : result2 = 100753;
		16'd7977 : result2 = 101227;
		16'd7978 : result2 = 101724;
		16'd7979 : result2 = 102243;
		16'd7980 : result2 = 102785;
		16'd7981 : result2 = 103350;
		16'd7982 : result2 = 103939;
		16'd7983 : result2 = 104552;
		16'd7984 : result2 = 105189;
		16'd7985 : result2 = 105851;
		16'd7986 : result2 = 106540;
		16'd8192 : result2 = 106066;
		16'd8193 : result2 = 104905;
		16'd8194 : result2 = 103812;
		16'd8195 : result2 = 102789;
		16'd8196 : result2 = 101838;
		16'd8197 : result2 = 100958;
		16'd8198 : result2 = 100147;
		16'd8199 : result2 = 99403;
		16'd8200 : result2 = 98725;
		16'd8201 : result2 = 98109;
		16'd8202 : result2 = 97553;
		16'd8203 : result2 = 97056;
		16'd8204 : result2 = 96613;
		16'd8205 : result2 = 96223;
		16'd8206 : result2 = 95884;
		16'd8207 : result2 = 95592;
		16'd8208 : result2 = 95347;
		16'd8209 : result2 = 95145;
		16'd8210 : result2 = 94985;
		16'd8211 : result2 = 94865;
		16'd8212 : result2 = 94783;
		16'd8213 : result2 = 94738;
		16'd8214 : result2 = 94728;
		16'd8215 : result2 = 94752;
		16'd8216 : result2 = 94809;
		16'd8217 : result2 = 94896;
		16'd8218 : result2 = 95014;
		16'd8219 : result2 = 95160;
		16'd8220 : result2 = 95335;
		16'd8221 : result2 = 95536;
		16'd8222 : result2 = 95764;
		16'd8223 : result2 = 96018;
		16'd8224 : result2 = 96297;
		16'd8225 : result2 = 96600;
		16'd8226 : result2 = 96927;
		16'd8227 : result2 = 97277;
		16'd8228 : result2 = 97651;
		16'd8229 : result2 = 98047;
		16'd8230 : result2 = 98466;
		16'd8231 : result2 = 98907;
		16'd8232 : result2 = 99370;
		16'd8233 : result2 = 99856;
		16'd8234 : result2 = 100363;
		16'd8235 : result2 = 100893;
		16'd8236 : result2 = 101446;
		16'd8237 : result2 = 102021;
		16'd8238 : result2 = 102619;
		16'd8239 : result2 = 103240;
		16'd8240 : result2 = 103886;
		16'd8241 : result2 = 104557;
		16'd8242 : result2 = 105253;
		16'd8448 : result2 = 104648;
		16'd8449 : result2 = 103399;
		16'd8450 : result2 = 102237;
		16'd8451 : result2 = 101161;
		16'd8452 : result2 = 100168;
		16'd8453 : result2 = 99256;
		16'd8454 : result2 = 98421;
		16'd8455 : result2 = 97661;
		16'd8456 : result2 = 96971;
		16'd8457 : result2 = 96349;
		16'd8458 : result2 = 95792;
		16'd8459 : result2 = 95295;
		16'd8460 : result2 = 94856;
		16'd8461 : result2 = 94472;
		16'd8462 : result2 = 94141;
		16'd8463 : result2 = 93859;
		16'd8464 : result2 = 93625;
		16'd8465 : result2 = 93435;
		16'd8466 : result2 = 93289;
		16'd8467 : result2 = 93183;
		16'd8468 : result2 = 93116;
		16'd8469 : result2 = 93086;
		16'd8470 : result2 = 93091;
		16'd8471 : result2 = 93130;
		16'd8472 : result2 = 93202;
		16'd8473 : result2 = 93305;
		16'd8474 : result2 = 93439;
		16'd8475 : result2 = 93601;
		16'd8476 : result2 = 93791;
		16'd8477 : result2 = 94008;
		16'd8478 : result2 = 94251;
		16'd8479 : result2 = 94520;
		16'd8480 : result2 = 94814;
		16'd8481 : result2 = 95131;
		16'd8482 : result2 = 95472;
		16'd8483 : result2 = 95837;
		16'd8484 : result2 = 96224;
		16'd8485 : result2 = 96633;
		16'd8486 : result2 = 97065;
		16'd8487 : result2 = 97519;
		16'd8488 : result2 = 97994;
		16'd8489 : result2 = 98492;
		16'd8490 : result2 = 99011;
		16'd8491 : result2 = 99552;
		16'd8492 : result2 = 100115;
		16'd8493 : result2 = 100700;
		16'd8494 : result2 = 101308;
		16'd8495 : result2 = 101939;
		16'd8496 : result2 = 102594;
		16'd8497 : result2 = 103272;
		16'd8498 : result2 = 103976;
		16'd8704 : result2 = 103121;
		16'd8705 : result2 = 101801;
		16'd8706 : result2 = 100583;
		16'd8707 : result2 = 99463;
		16'd8708 : result2 = 98438;
		16'd8709 : result2 = 97501;
		16'd8710 : result2 = 96649;
		16'd8711 : result2 = 95877;
		16'd8712 : result2 = 95181;
		16'd8713 : result2 = 94557;
		16'd8714 : result2 = 94001;
		16'd8715 : result2 = 93508;
		16'd8716 : result2 = 93076;
		16'd8717 : result2 = 92701;
		16'd8718 : result2 = 92380;
		16'd8719 : result2 = 92111;
		16'd8720 : result2 = 91890;
		16'd8721 : result2 = 91714;
		16'd8722 : result2 = 91582;
		16'd8723 : result2 = 91492;
		16'd8724 : result2 = 91441;
		16'd8725 : result2 = 91427;
		16'd8726 : result2 = 91449;
		16'd8727 : result2 = 91505;
		16'd8728 : result2 = 91593;
		16'd8729 : result2 = 91713;
		16'd8730 : result2 = 91863;
		16'd8731 : result2 = 92042;
		16'd8732 : result2 = 92248;
		16'd8733 : result2 = 92481;
		16'd8734 : result2 = 92740;
		16'd8735 : result2 = 93025;
		16'd8736 : result2 = 93334;
		16'd8737 : result2 = 93666;
		16'd8738 : result2 = 94022;
		16'd8739 : result2 = 94401;
		16'd8740 : result2 = 94802;
		16'd8741 : result2 = 95226;
		16'd8742 : result2 = 95671;
		16'd8743 : result2 = 96138;
		16'd8744 : result2 = 96626;
		16'd8745 : result2 = 97135;
		16'd8746 : result2 = 97666;
		16'd8747 : result2 = 98219;
		16'd8748 : result2 = 98793;
		16'd8749 : result2 = 99389;
		16'd8750 : result2 = 100007;
		16'd8751 : result2 = 100647;
		16'd8752 : result2 = 101311;
		16'd8753 : result2 = 101999;
		16'd8754 : result2 = 102711;
		16'd8960 : result2 = 101483;
		16'd8961 : result2 = 100107;
		16'd8962 : result2 = 98847;
		16'd8963 : result2 = 97694;
		16'd8964 : result2 = 96644;
		16'd8965 : result2 = 95691;
		16'd8966 : result2 = 94828;
		16'd8967 : result2 = 94050;
		16'd8968 : result2 = 93353;
		16'd8969 : result2 = 92731;
		16'd8970 : result2 = 92179;
		16'd8971 : result2 = 91695;
		16'd8972 : result2 = 91273;
		16'd8973 : result2 = 90910;
		16'd8974 : result2 = 90602;
		16'd8975 : result2 = 90347;
		16'd8976 : result2 = 90141;
		16'd8977 : result2 = 89981;
		16'd8978 : result2 = 89866;
		16'd8979 : result2 = 89793;
		16'd8980 : result2 = 89759;
		16'd8981 : result2 = 89763;
		16'd8982 : result2 = 89802;
		16'd8983 : result2 = 89876;
		16'd8984 : result2 = 89982;
		16'd8985 : result2 = 90120;
		16'd8986 : result2 = 90287;
		16'd8987 : result2 = 90483;
		16'd8988 : result2 = 90706;
		16'd8989 : result2 = 90956;
		16'd8990 : result2 = 91232;
		16'd8991 : result2 = 91533;
		16'd8992 : result2 = 91858;
		16'd8993 : result2 = 92206;
		16'd8994 : result2 = 92577;
		16'd8995 : result2 = 92971;
		16'd8996 : result2 = 93387;
		16'd8997 : result2 = 93824;
		16'd8998 : result2 = 94283;
		16'd8999 : result2 = 94763;
		16'd9000 : result2 = 95264;
		16'd9001 : result2 = 95787;
		16'd9002 : result2 = 96330;
		16'd9003 : result2 = 96894;
		16'd9004 : result2 = 97479;
		16'd9005 : result2 = 98086;
		16'd9006 : result2 = 98715;
		16'd9007 : result2 = 99366;
		16'd9008 : result2 = 100039;
		16'd9009 : result2 = 100736;
		16'd9010 : result2 = 101457;
		16'd9216 : result2 = 99733;
		16'd9217 : result2 = 98318;
		16'd9218 : result2 = 97027;
		16'd9219 : result2 = 95852;
		16'd9220 : result2 = 94787;
		16'd9221 : result2 = 93824;
		16'd9222 : result2 = 92957;
		16'd9223 : result2 = 92179;
		16'd9224 : result2 = 91485;
		16'd9225 : result2 = 90870;
		16'd9226 : result2 = 90328;
		16'd9227 : result2 = 89855;
		16'd9228 : result2 = 89446;
		16'd9229 : result2 = 89097;
		16'd9230 : result2 = 88805;
		16'd9231 : result2 = 88567;
		16'd9232 : result2 = 88378;
		16'd9233 : result2 = 88237;
		16'd9234 : result2 = 88140;
		16'd9235 : result2 = 88085;
		16'd9236 : result2 = 88070;
		16'd9237 : result2 = 88093;
		16'd9238 : result2 = 88152;
		16'd9239 : result2 = 88244;
		16'd9240 : result2 = 88369;
		16'd9241 : result2 = 88525;
		16'd9242 : result2 = 88711;
		16'd9243 : result2 = 88925;
		16'd9244 : result2 = 89166;
		16'd9245 : result2 = 89434;
		16'd9246 : result2 = 89727;
		16'd9247 : result2 = 90045;
		16'd9248 : result2 = 90386;
		16'd9249 : result2 = 90750;
		16'd9250 : result2 = 91137;
		16'd9251 : result2 = 91547;
		16'd9252 : result2 = 91977;
		16'd9253 : result2 = 92429;
		16'd9254 : result2 = 92903;
		16'd9255 : result2 = 93397;
		16'd9256 : result2 = 93911;
		16'd9257 : result2 = 94446;
		16'd9258 : result2 = 95002;
		16'd9259 : result2 = 95578;
		16'd9260 : result2 = 96176;
		16'd9261 : result2 = 96794;
		16'd9262 : result2 = 97433;
		16'd9263 : result2 = 98094;
		16'd9264 : result2 = 98778;
		16'd9265 : result2 = 99484;
		16'd9266 : result2 = 100214;
		16'd9472 : result2 = 97874;
		16'd9473 : result2 = 96432;
		16'd9474 : result2 = 95123;
		16'd9475 : result2 = 93936;
		16'd9476 : result2 = 92864;
		16'd9477 : result2 = 91900;
		16'd9478 : result2 = 91035;
		16'd9479 : result2 = 90263;
		16'd9480 : result2 = 89578;
		16'd9481 : result2 = 88974;
		16'd9482 : result2 = 88446;
		16'd9483 : result2 = 87987;
		16'd9484 : result2 = 87595;
		16'd9485 : result2 = 87264;
		16'd9486 : result2 = 86991;
		16'd9487 : result2 = 86771;
		16'd9488 : result2 = 86602;
		16'd9489 : result2 = 86481;
		16'd9490 : result2 = 86405;
		16'd9491 : result2 = 86370;
		16'd9492 : result2 = 86376;
		16'd9493 : result2 = 86419;
		16'd9494 : result2 = 86498;
		16'd9495 : result2 = 86610;
		16'd9496 : result2 = 86755;
		16'd9497 : result2 = 86931;
		16'd9498 : result2 = 87136;
		16'd9499 : result2 = 87369;
		16'd9500 : result2 = 87629;
		16'd9501 : result2 = 87914;
		16'd9502 : result2 = 88225;
		16'd9503 : result2 = 88560;
		16'd9504 : result2 = 88919;
		16'd9505 : result2 = 89300;
		16'd9506 : result2 = 89703;
		16'd9507 : result2 = 90128;
		16'd9508 : result2 = 90574;
		16'd9509 : result2 = 91042;
		16'd9510 : result2 = 91529;
		16'd9511 : result2 = 92037;
		16'd9512 : result2 = 92566;
		16'd9513 : result2 = 93114;
		16'd9514 : result2 = 93683;
		16'd9515 : result2 = 94272;
		16'd9516 : result2 = 94881;
		16'd9517 : result2 = 95511;
		16'd9518 : result2 = 96162;
		16'd9519 : result2 = 96833;
		16'd9520 : result2 = 97527;
		16'd9521 : result2 = 98243;
		16'd9522 : result2 = 98983;
		16'd9728 : result2 = 95906;
		16'd9729 : result2 = 94451;
		16'd9730 : result2 = 93135;
		16'd9731 : result2 = 91946;
		16'd9732 : result2 = 90876;
		16'd9733 : result2 = 89918;
		16'd9734 : result2 = 89062;
		16'd9735 : result2 = 88303;
		16'd9736 : result2 = 87632;
		16'd9737 : result2 = 87044;
		16'd9738 : result2 = 86533;
		16'd9739 : result2 = 86094;
		16'd9740 : result2 = 85721;
		16'd9741 : result2 = 85411;
		16'd9742 : result2 = 85159;
		16'd9743 : result2 = 84961;
		16'd9744 : result2 = 84814;
		16'd9745 : result2 = 84715;
		16'd9746 : result2 = 84660;
		16'd9747 : result2 = 84648;
		16'd9748 : result2 = 84675;
		16'd9749 : result2 = 84740;
		16'd9750 : result2 = 84841;
		16'd9751 : result2 = 84974;
		16'd9752 : result2 = 85140;
		16'd9753 : result2 = 85336;
		16'd9754 : result2 = 85561;
		16'd9755 : result2 = 85814;
		16'd9756 : result2 = 86093;
		16'd9757 : result2 = 86398;
		16'd9758 : result2 = 86728;
		16'd9759 : result2 = 87081;
		16'd9760 : result2 = 87457;
		16'd9761 : result2 = 87855;
		16'd9762 : result2 = 88275;
		16'd9763 : result2 = 88716;
		16'd9764 : result2 = 89179;
		16'd9765 : result2 = 89661;
		16'd9766 : result2 = 90164;
		16'd9767 : result2 = 90686;
		16'd9768 : result2 = 91229;
		16'd9769 : result2 = 91791;
		16'd9770 : result2 = 92373;
		16'd9771 : result2 = 92975;
		16'd9772 : result2 = 93596;
		16'd9773 : result2 = 94238;
		16'd9774 : result2 = 94900;
		16'd9775 : result2 = 95583;
		16'd9776 : result2 = 96287;
		16'd9777 : result2 = 97014;
		16'd9778 : result2 = 97763;
		16'd9984 : result2 = 93831;
		16'd9985 : result2 = 92376;
		16'd9986 : result2 = 91064;
		16'd9987 : result2 = 89882;
		16'd9988 : result2 = 88824;
		16'd9989 : result2 = 87879;
		16'd9990 : result2 = 87039;
		16'd9991 : result2 = 86297;
		16'd9992 : result2 = 85646;
		16'd9993 : result2 = 85079;
		16'd9994 : result2 = 84590;
		16'd9995 : result2 = 84174;
		16'd9996 : result2 = 83824;
		16'd9997 : result2 = 83538;
		16'd9998 : result2 = 83310;
		16'd9999 : result2 = 83136;
		16'd10000 : result2 = 83014;
		16'd10001 : result2 = 82939;
		16'd10002 : result2 = 82908;
		16'd10003 : result2 = 82919;
		16'd10004 : result2 = 82970;
		16'd10005 : result2 = 83058;
		16'd10006 : result2 = 83181;
		16'd10007 : result2 = 83337;
		16'd10008 : result2 = 83525;
		16'd10009 : result2 = 83743;
		16'd10010 : result2 = 83989;
		16'd10011 : result2 = 84262;
		16'd10012 : result2 = 84561;
		16'd10013 : result2 = 84886;
		16'd10014 : result2 = 85234;
		16'd10015 : result2 = 85606;
		16'd10016 : result2 = 86000;
		16'd10017 : result2 = 86416;
		16'd10018 : result2 = 86853;
		16'd10019 : result2 = 87312;
		16'd10020 : result2 = 87790;
		16'd10021 : result2 = 88288;
		16'd10022 : result2 = 88806;
		16'd10023 : result2 = 89344;
		16'd10024 : result2 = 89901;
		16'd10025 : result2 = 90477;
		16'd10026 : result2 = 91072;
		16'd10027 : result2 = 91687;
		16'd10028 : result2 = 92321;
		16'd10029 : result2 = 92975;
		16'd10030 : result2 = 93649;
		16'd10031 : result2 = 94343;
		16'd10032 : result2 = 95058;
		16'd10033 : result2 = 95795;
		16'd10034 : result2 = 96554;
		16'd10240 : result2 = 91652;
		16'd10241 : result2 = 90209;
		16'd10242 : result2 = 88910;
		16'd10243 : result2 = 87746;
		16'd10244 : result2 = 86707;
		16'd10245 : result2 = 85783;
		16'd10246 : result2 = 84966;
		16'd10247 : result2 = 84248;
		16'd10248 : result2 = 83622;
		16'd10249 : result2 = 83081;
		16'd10250 : result2 = 82618;
		16'd10251 : result2 = 82228;
		16'd10252 : result2 = 81906;
		16'd10253 : result2 = 81646;
		16'd10254 : result2 = 81445;
		16'd10255 : result2 = 81298;
		16'd10256 : result2 = 81202;
		16'd10257 : result2 = 81153;
		16'd10258 : result2 = 81148;
		16'd10259 : result2 = 81185;
		16'd10260 : result2 = 81261;
		16'd10261 : result2 = 81373;
		16'd10262 : result2 = 81520;
		16'd10263 : result2 = 81700;
		16'd10264 : result2 = 81910;
		16'd10265 : result2 = 82150;
		16'd10266 : result2 = 82418;
		16'd10267 : result2 = 82713;
		16'd10268 : result2 = 83033;
		16'd10269 : result2 = 83378;
		16'd10270 : result2 = 83746;
		16'd10271 : result2 = 84137;
		16'd10272 : result2 = 84550;
		16'd10273 : result2 = 84984;
		16'd10274 : result2 = 85439;
		16'd10275 : result2 = 85914;
		16'd10276 : result2 = 86409;
		16'd10277 : result2 = 86924;
		16'd10278 : result2 = 87457;
		16'd10279 : result2 = 88010;
		16'd10280 : result2 = 88582;
		16'd10281 : result2 = 89172;
		16'd10282 : result2 = 89781;
		16'd10283 : result2 = 90409;
		16'd10284 : result2 = 91056;
		16'd10285 : result2 = 91723;
		16'd10286 : result2 = 92409;
		16'd10287 : result2 = 93115;
		16'd10288 : result2 = 93841;
		16'd10289 : result2 = 94588;
		16'd10290 : result2 = 95357;
		16'd10496 : result2 = 89371;
		16'd10497 : result2 = 87951;
		16'd10498 : result2 = 86677;
		16'd10499 : result2 = 85539;
		16'd10500 : result2 = 84527;
		16'd10501 : result2 = 83632;
		16'd10502 : result2 = 82844;
		16'd10503 : result2 = 82156;
		16'd10504 : result2 = 81560;
		16'd10505 : result2 = 81050;
		16'd10506 : result2 = 80618;
		16'd10507 : result2 = 80258;
		16'd10508 : result2 = 79967;
		16'd10509 : result2 = 79737;
		16'd10510 : result2 = 79565;
		16'd10511 : result2 = 79448;
		16'd10512 : result2 = 79380;
		16'd10513 : result2 = 79359;
		16'd10514 : result2 = 79382;
		16'd10515 : result2 = 79446;
		16'd10516 : result2 = 79548;
		16'd10517 : result2 = 79686;
		16'd10518 : result2 = 79858;
		16'd10519 : result2 = 80063;
		16'd10520 : result2 = 80297;
		16'd10521 : result2 = 80560;
		16'd10522 : result2 = 80851;
		16'd10523 : result2 = 81168;
		16'd10524 : result2 = 81509;
		16'd10525 : result2 = 81875;
		16'd10526 : result2 = 82263;
		16'd10527 : result2 = 82674;
		16'd10528 : result2 = 83106;
		16'd10529 : result2 = 83559;
		16'd10530 : result2 = 84032;
		16'd10531 : result2 = 84524;
		16'd10532 : result2 = 85036;
		16'd10533 : result2 = 85567;
		16'd10534 : result2 = 86117;
		16'd10535 : result2 = 86685;
		16'd10536 : result2 = 87272;
		16'd10537 : result2 = 87877;
		16'd10538 : result2 = 88500;
		16'd10539 : result2 = 89142;
		16'd10540 : result2 = 89802;
		16'd10541 : result2 = 90481;
		16'd10542 : result2 = 91179;
		16'd10543 : result2 = 91897;
		16'd10544 : result2 = 92635;
		16'd10545 : result2 = 93393;
		16'd10546 : result2 = 94172;
		16'd10752 : result2 = 86992;
		16'd10753 : result2 = 85605;
		16'd10754 : result2 = 84366;
		16'd10755 : result2 = 83263;
		16'd10756 : result2 = 82286;
		16'd10757 : result2 = 81427;
		16'd10758 : result2 = 80675;
		16'd10759 : result2 = 80023;
		16'd10760 : result2 = 79463;
		16'd10761 : result2 = 78988;
		16'd10762 : result2 = 78591;
		16'd10763 : result2 = 78266;
		16'd10764 : result2 = 78008;
		16'd10765 : result2 = 77811;
		16'd10766 : result2 = 77672;
		16'd10767 : result2 = 77586;
		16'd10768 : result2 = 77549;
		16'd10769 : result2 = 77559;
		16'd10770 : result2 = 77611;
		16'd10771 : result2 = 77703;
		16'd10772 : result2 = 77833;
		16'd10773 : result2 = 77998;
		16'd10774 : result2 = 78197;
		16'd10775 : result2 = 78427;
		16'd10776 : result2 = 78686;
		16'd10777 : result2 = 78973;
		16'd10778 : result2 = 79287;
		16'd10779 : result2 = 79627;
		16'd10780 : result2 = 79991;
		16'd10781 : result2 = 80378;
		16'd10782 : result2 = 80787;
		16'd10783 : result2 = 81218;
		16'd10784 : result2 = 81669;
		16'd10785 : result2 = 82141;
		16'd10786 : result2 = 82633;
		16'd10787 : result2 = 83143;
		16'd10788 : result2 = 83673;
		16'd10789 : result2 = 84220;
		16'd10790 : result2 = 84786;
		16'd10791 : result2 = 85370;
		16'd10792 : result2 = 85972;
		16'd10793 : result2 = 86592;
		16'd10794 : result2 = 87230;
		16'd10795 : result2 = 87885;
		16'd10796 : result2 = 88559;
		16'd10797 : result2 = 89251;
		16'd10798 : result2 = 89961;
		16'd10799 : result2 = 90691;
		16'd10800 : result2 = 91440;
		16'd10801 : result2 = 92209;
		16'd10802 : result2 = 93000;
		16'd11008 : result2 = 84517;
		16'd11009 : result2 = 83174;
		16'd11010 : result2 = 81979;
		16'd11011 : result2 = 80920;
		16'd11012 : result2 = 79987;
		16'd11013 : result2 = 79171;
		16'd11014 : result2 = 78462;
		16'd11015 : result2 = 77851;
		16'd11016 : result2 = 77332;
		16'd11017 : result2 = 76897;
		16'd11018 : result2 = 76539;
		16'd11019 : result2 = 76252;
		16'd11020 : result2 = 76031;
		16'd11021 : result2 = 75870;
		16'd11022 : result2 = 75766;
		16'd11023 : result2 = 75714;
		16'd11024 : result2 = 75711;
		16'd11025 : result2 = 75752;
		16'd11026 : result2 = 75835;
		16'd11027 : result2 = 75958;
		16'd11028 : result2 = 76117;
		16'd11029 : result2 = 76310;
		16'd11030 : result2 = 76536;
		16'd11031 : result2 = 76793;
		16'd11032 : result2 = 77078;
		16'd11033 : result2 = 77390;
		16'd11034 : result2 = 77728;
		16'd11035 : result2 = 78091;
		16'd11036 : result2 = 78478;
		16'd11037 : result2 = 78887;
		16'd11038 : result2 = 79317;
		16'd11039 : result2 = 79769;
		16'd11040 : result2 = 80241;
		16'd11041 : result2 = 80732;
		16'd11042 : result2 = 81242;
		16'd11043 : result2 = 81771;
		16'd11044 : result2 = 82318;
		16'd11045 : result2 = 82883;
		16'd11046 : result2 = 83465;
		16'd11047 : result2 = 84065;
		16'd11048 : result2 = 84683;
		16'd11049 : result2 = 85317;
		16'd11050 : result2 = 85970;
		16'd11051 : result2 = 86639;
		16'd11052 : result2 = 87326;
		16'd11053 : result2 = 88031;
		16'd11054 : result2 = 88755;
		16'd11055 : result2 = 89496;
		16'd11056 : result2 = 90257;
		16'd11057 : result2 = 91038;
		16'd11058 : result2 = 91839;
		16'd11264 : result2 = 81949;
		16'd11265 : result2 = 80661;
		16'd11266 : result2 = 79519;
		16'd11267 : result2 = 78513;
		16'd11268 : result2 = 77632;
		16'd11269 : result2 = 76866;
		16'd11270 : result2 = 76205;
		16'd11271 : result2 = 75643;
		16'd11272 : result2 = 75170;
		16'd11273 : result2 = 74779;
		16'd11274 : result2 = 74464;
		16'd11275 : result2 = 74219;
		16'd11276 : result2 = 74038;
		16'd11277 : result2 = 73916;
		16'd11278 : result2 = 73850;
		16'd11279 : result2 = 73834;
		16'd11280 : result2 = 73866;
		16'd11281 : result2 = 73941;
		16'd11282 : result2 = 74057;
		16'd11283 : result2 = 74211;
		16'd11284 : result2 = 74401;
		16'd11285 : result2 = 74624;
		16'd11286 : result2 = 74878;
		16'd11287 : result2 = 75162;
		16'd11288 : result2 = 75474;
		16'd11289 : result2 = 75812;
		16'd11290 : result2 = 76175;
		16'd11291 : result2 = 76562;
		16'd11292 : result2 = 76972;
		16'd11293 : result2 = 77403;
		16'd11294 : result2 = 77856;
		16'd11295 : result2 = 78328;
		16'd11296 : result2 = 78820;
		16'd11297 : result2 = 79331;
		16'd11298 : result2 = 79861;
		16'd11299 : result2 = 80408;
		16'd11300 : result2 = 80973;
		16'd11301 : result2 = 81555;
		16'd11302 : result2 = 82154;
		16'd11303 : result2 = 82771;
		16'd11304 : result2 = 83404;
		16'd11305 : result2 = 84054;
		16'd11306 : result2 = 84721;
		16'd11307 : result2 = 85404;
		16'd11308 : result2 = 86105;
		16'd11309 : result2 = 86824;
		16'd11310 : result2 = 87560;
		16'd11311 : result2 = 88314;
		16'd11312 : result2 = 89087;
		16'd11313 : result2 = 89879;
		16'd11314 : result2 = 90691;
		16'd11520 : result2 = 79294;
		16'd11521 : result2 = 78070;
		16'd11522 : result2 = 76992;
		16'd11523 : result2 = 76047;
		16'd11524 : result2 = 75224;
		16'd11525 : result2 = 74515;
		16'd11526 : result2 = 73910;
		16'd11527 : result2 = 73400;
		16'd11528 : result2 = 72978;
		16'd11529 : result2 = 72636;
		16'd11530 : result2 = 72368;
		16'd11531 : result2 = 72168;
		16'd11532 : result2 = 72031;
		16'd11533 : result2 = 71951;
		16'd11534 : result2 = 71925;
		16'd11535 : result2 = 71947;
		16'd11536 : result2 = 72016;
		16'd11537 : result2 = 72127;
		16'd11538 : result2 = 72277;
		16'd11539 : result2 = 72464;
		16'd11540 : result2 = 72686;
		16'd11541 : result2 = 72939;
		16'd11542 : result2 = 73223;
		16'd11543 : result2 = 73536;
		16'd11544 : result2 = 73875;
		16'd11545 : result2 = 74239;
		16'd11546 : result2 = 74628;
		16'd11547 : result2 = 75040;
		16'd11548 : result2 = 75473;
		16'd11549 : result2 = 75928;
		16'd11550 : result2 = 76402;
		16'd11551 : result2 = 76896;
		16'd11552 : result2 = 77409;
		16'd11553 : result2 = 77940;
		16'd11554 : result2 = 78489;
		16'd11555 : result2 = 79055;
		16'd11556 : result2 = 79638;
		16'd11557 : result2 = 80238;
		16'd11558 : result2 = 80854;
		16'd11559 : result2 = 81487;
		16'd11560 : result2 = 82136;
		16'd11561 : result2 = 82801;
		16'd11562 : result2 = 83483;
		16'd11563 : result2 = 84181;
		16'd11564 : result2 = 84896;
		16'd11565 : result2 = 85628;
		16'd11566 : result2 = 86377;
		16'd11567 : result2 = 87144;
		16'd11568 : result2 = 87929;
		16'd11569 : result2 = 88733;
		16'd11570 : result2 = 89556;
		16'd11776 : result2 = 76555;
		16'd11777 : result2 = 75406;
		16'd11778 : result2 = 74400;
		16'd11779 : result2 = 73524;
		16'd11780 : result2 = 72769;
		16'd11781 : result2 = 72123;
		16'd11782 : result2 = 71579;
		16'd11783 : result2 = 71128;
		16'd11784 : result2 = 70761;
		16'd11785 : result2 = 70472;
		16'd11786 : result2 = 70255;
		16'd11787 : result2 = 70104;
		16'd11788 : result2 = 70012;
		16'd11789 : result2 = 69977;
		16'd11790 : result2 = 69993;
		16'd11791 : result2 = 70056;
		16'd11792 : result2 = 70164;
		16'd11793 : result2 = 70312;
		16'd11794 : result2 = 70498;
		16'd11795 : result2 = 70719;
		16'd11796 : result2 = 70973;
		16'd11797 : result2 = 71259;
		16'd11798 : result2 = 71573;
		16'd11799 : result2 = 71914;
		16'd11800 : result2 = 72282;
		16'd11801 : result2 = 72673;
		16'd11802 : result2 = 73088;
		16'd11803 : result2 = 73525;
		16'd11804 : result2 = 73983;
		16'd11805 : result2 = 74461;
		16'd11806 : result2 = 74958;
		16'd11807 : result2 = 75474;
		16'd11808 : result2 = 76008;
		16'd11809 : result2 = 76559;
		16'd11810 : result2 = 77128;
		16'd11811 : result2 = 77713;
		16'd11812 : result2 = 78314;
		16'd11813 : result2 = 78932;
		16'd11814 : result2 = 79565;
		16'd11815 : result2 = 80215;
		16'd11816 : result2 = 80880;
		16'd11817 : result2 = 81561;
		16'd11818 : result2 = 82258;
		16'd11819 : result2 = 82970;
		16'd11820 : result2 = 83699;
		16'd11821 : result2 = 84445;
		16'd11822 : result2 = 85207;
		16'd11823 : result2 = 85987;
		16'd11824 : result2 = 86784;
		16'd11825 : result2 = 87600;
		16'd11826 : result2 = 88435;
		16'd12032 : result2 = 73738;
		16'd12033 : result2 = 72675;
		16'd12034 : result2 = 71749;
		16'd12035 : result2 = 70951;
		16'd12036 : result2 = 70269;
		16'd12037 : result2 = 69694;
		16'd12038 : result2 = 69216;
		16'd12039 : result2 = 68828;
		16'd12040 : result2 = 68522;
		16'd12041 : result2 = 68290;
		16'd12042 : result2 = 68127;
		16'd12043 : result2 = 68027;
		16'd12044 : result2 = 67985;
		16'd12045 : result2 = 67996;
		16'd12046 : result2 = 68057;
		16'd12047 : result2 = 68162;
		16'd12048 : result2 = 68310;
		16'd12049 : result2 = 68497;
		16'd12050 : result2 = 68720;
		16'd12051 : result2 = 68977;
		16'd12052 : result2 = 69265;
		16'd12053 : result2 = 69583;
		16'd12054 : result2 = 69928;
		16'd12055 : result2 = 70300;
		16'd12056 : result2 = 70696;
		16'd12057 : result2 = 71115;
		16'd12058 : result2 = 71557;
		16'd12059 : result2 = 72019;
		16'd12060 : result2 = 72502;
		16'd12061 : result2 = 73003;
		16'd12062 : result2 = 73524;
		16'd12063 : result2 = 74062;
		16'd12064 : result2 = 74617;
		16'd12065 : result2 = 75189;
		16'd12066 : result2 = 75777;
		16'd12067 : result2 = 76382;
		16'd12068 : result2 = 77002;
		16'd12069 : result2 = 77637;
		16'd12070 : result2 = 78288;
		16'd12071 : result2 = 78954;
		16'd12072 : result2 = 79636;
		16'd12073 : result2 = 80332;
		16'd12074 : result2 = 81044;
		16'd12075 : result2 = 81772;
		16'd12076 : result2 = 82515;
		16'd12077 : result2 = 83274;
		16'd12078 : result2 = 84050;
		16'd12079 : result2 = 84842;
		16'd12080 : result2 = 85652;
		16'd12081 : result2 = 86479;
		16'd12082 : result2 = 87326;
		16'd12288 : result2 = 70850;
		16'd12289 : result2 = 69881;
		16'd12290 : result2 = 69046;
		16'd12291 : result2 = 68333;
		16'd12292 : result2 = 67731;
		16'd12293 : result2 = 67232;
		16'd12294 : result2 = 66827;
		16'd12295 : result2 = 66506;
		16'd12296 : result2 = 66264;
		16'd12297 : result2 = 66093;
		16'd12298 : result2 = 65987;
		16'd12299 : result2 = 65942;
		16'd12300 : result2 = 65951;
		16'd12301 : result2 = 66011;
		16'd12302 : result2 = 66118;
		16'd12303 : result2 = 66268;
		16'd12304 : result2 = 66458;
		16'd12305 : result2 = 66685;
		16'd12306 : result2 = 66946;
		16'd12307 : result2 = 67240;
		16'd12308 : result2 = 67563;
		16'd12309 : result2 = 67914;
		16'd12310 : result2 = 68291;
		16'd12311 : result2 = 68693;
		16'd12312 : result2 = 69119;
		16'd12313 : result2 = 69566;
		16'd12314 : result2 = 70035;
		16'd12315 : result2 = 70523;
		16'd12316 : result2 = 71031;
		16'd12317 : result2 = 71557;
		16'd12318 : result2 = 72100;
		16'd12319 : result2 = 72660;
		16'd12320 : result2 = 73237;
		16'd12321 : result2 = 73830;
		16'd12322 : result2 = 74439;
		16'd12323 : result2 = 75062;
		16'd12324 : result2 = 75701;
		16'd12325 : result2 = 76355;
		16'd12326 : result2 = 77023;
		16'd12327 : result2 = 77706;
		16'd12328 : result2 = 78404;
		16'd12329 : result2 = 79116;
		16'd12330 : result2 = 79844;
		16'd12331 : result2 = 80586;
		16'd12332 : result2 = 81343;
		16'd12333 : result2 = 82116;
		16'd12334 : result2 = 82905;
		16'd12335 : result2 = 83711;
		16'd12336 : result2 = 84533;
		16'd12337 : result2 = 85373;
		16'd12338 : result2 = 86231;
		16'd12544 : result2 = 67898;
		16'd12545 : result2 = 67033;
		16'd12546 : result2 = 66296;
		16'd12547 : result2 = 65675;
		16'd12548 : result2 = 65161;
		16'd12549 : result2 = 64744;
		16'd12550 : result2 = 64415;
		16'd12551 : result2 = 64167;
		16'd12552 : result2 = 63992;
		16'd12553 : result2 = 63885;
		16'd12554 : result2 = 63840;
		16'd12555 : result2 = 63851;
		16'd12556 : result2 = 63915;
		16'd12557 : result2 = 64026;
		16'd12558 : result2 = 64181;
		16'd12559 : result2 = 64376;
		16'd12560 : result2 = 64609;
		16'd12561 : result2 = 64878;
		16'd12562 : result2 = 65178;
		16'd12563 : result2 = 65509;
		16'd12564 : result2 = 65868;
		16'd12565 : result2 = 66253;
		16'd12566 : result2 = 66663;
		16'd12567 : result2 = 67096;
		16'd12568 : result2 = 67551;
		16'd12569 : result2 = 68028;
		16'd12570 : result2 = 68524;
		16'd12571 : result2 = 69038;
		16'd12572 : result2 = 69571;
		16'd12573 : result2 = 70121;
		16'd12574 : result2 = 70688;
		16'd12575 : result2 = 71271;
		16'd12576 : result2 = 71870;
		16'd12577 : result2 = 72484;
		16'd12578 : result2 = 73112;
		16'd12579 : result2 = 73756;
		16'd12580 : result2 = 74413;
		16'd12581 : result2 = 75085;
		16'd12582 : result2 = 75771;
		16'd12583 : result2 = 76471;
		16'd12584 : result2 = 77185;
		16'd12585 : result2 = 77913;
		16'd12586 : result2 = 78656;
		16'd12587 : result2 = 79413;
		16'd12588 : result2 = 80185;
		16'd12589 : result2 = 80972;
		16'd12590 : result2 = 81774;
		16'd12591 : result2 = 82593;
		16'd12592 : result2 = 83427;
		16'd12593 : result2 = 84280;
		16'd12594 : result2 = 85150;
		16'd12800 : result2 = 64891;
		16'd12801 : result2 = 64139;
		16'd12802 : result2 = 63508;
		16'd12803 : result2 = 62986;
		16'd12804 : result2 = 62565;
		16'd12805 : result2 = 62234;
		16'd12806 : result2 = 61986;
		16'd12807 : result2 = 61814;
		16'd12808 : result2 = 61711;
		16'd12809 : result2 = 61671;
		16'd12810 : result2 = 61688;
		16'd12811 : result2 = 61759;
		16'd12812 : result2 = 61878;
		16'd12813 : result2 = 62041;
		16'd12814 : result2 = 62246;
		16'd12815 : result2 = 62489;
		16'd12816 : result2 = 62766;
		16'd12817 : result2 = 63077;
		16'd12818 : result2 = 63417;
		16'd12819 : result2 = 63786;
		16'd12820 : result2 = 64181;
		16'd12821 : result2 = 64601;
		16'd12822 : result2 = 65044;
		16'd12823 : result2 = 65509;
		16'd12824 : result2 = 65995;
		16'd12825 : result2 = 66500;
		16'd12826 : result2 = 67024;
		16'd12827 : result2 = 67565;
		16'd12828 : result2 = 68124;
		16'd12829 : result2 = 68698;
		16'd12830 : result2 = 69289;
		16'd12831 : result2 = 69895;
		16'd12832 : result2 = 70515;
		16'd12833 : result2 = 71150;
		16'd12834 : result2 = 71799;
		16'd12835 : result2 = 72462;
		16'd12836 : result2 = 73138;
		16'd12837 : result2 = 73828;
		16'd12838 : result2 = 74532;
		16'd12839 : result2 = 75249;
		16'd12840 : result2 = 75980;
		16'd12841 : result2 = 76724;
		16'd12842 : result2 = 77482;
		16'd12843 : result2 = 78254;
		16'd12844 : result2 = 79040;
		16'd12845 : result2 = 79841;
		16'd12846 : result2 = 80657;
		16'd12847 : result2 = 81489;
		16'd12848 : result2 = 82336;
		16'd12849 : result2 = 83201;
		16'd12850 : result2 = 84082;
		16'd13056 : result2 = 61840;
		16'd13057 : result2 = 61209;
		16'd13058 : result2 = 60690;
		16'd13059 : result2 = 60273;
		16'd13060 : result2 = 59949;
		16'd13061 : result2 = 59710;
		16'd13062 : result2 = 59547;
		16'd13063 : result2 = 59454;
		16'd13064 : result2 = 59425;
		16'd13065 : result2 = 59454;
		16'd13066 : result2 = 59537;
		16'd13067 : result2 = 59668;
		16'd13068 : result2 = 59844;
		16'd13069 : result2 = 60062;
		16'd13070 : result2 = 60318;
		16'd13071 : result2 = 60608;
		16'd13072 : result2 = 60931;
		16'd13073 : result2 = 61285;
		16'd13074 : result2 = 61666;
		16'd13075 : result2 = 62074;
		16'd13076 : result2 = 62506;
		16'd13077 : result2 = 62961;
		16'd13078 : result2 = 63438;
		16'd13079 : result2 = 63935;
		16'd13080 : result2 = 64451;
		16'd13081 : result2 = 64985;
		16'd13082 : result2 = 65537;
		16'd13083 : result2 = 66105;
		16'd13084 : result2 = 66689;
		16'd13085 : result2 = 67289;
		16'd13086 : result2 = 67903;
		16'd13087 : result2 = 68531;
		16'd13088 : result2 = 69174;
		16'd13089 : result2 = 69830;
		16'd13090 : result2 = 70499;
		16'd13091 : result2 = 71182;
		16'd13092 : result2 = 71877;
		16'd13093 : result2 = 72586;
		16'd13094 : result2 = 73307;
		16'd13095 : result2 = 74041;
		16'd13096 : result2 = 74788;
		16'd13097 : result2 = 75549;
		16'd13098 : result2 = 76322;
		16'd13099 : result2 = 77109;
		16'd13100 : result2 = 77910;
		16'd13101 : result2 = 78725;
		16'd13102 : result2 = 79554;
		16'd13103 : result2 = 80399;
		16'd13104 : result2 = 81259;
		16'd13105 : result2 = 82136;
		16'd13106 : result2 = 83030;
		16'd13312 : result2 = 58754;
		16'd13313 : result2 = 58251;
		16'd13314 : result2 = 57851;
		16'd13315 : result2 = 57544;
		16'd13316 : result2 = 57323;
		16'd13317 : result2 = 57178;
		16'd13318 : result2 = 57103;
		16'd13319 : result2 = 57092;
		16'd13320 : result2 = 57140;
		16'd13321 : result2 = 57240;
		16'd13322 : result2 = 57389;
		16'd13323 : result2 = 57583;
		16'd13324 : result2 = 57818;
		16'd13325 : result2 = 58091;
		16'd13326 : result2 = 58398;
		16'd13327 : result2 = 58738;
		16'd13328 : result2 = 59107;
		16'd13329 : result2 = 59504;
		16'd13330 : result2 = 59927;
		16'd13331 : result2 = 60374;
		16'd13332 : result2 = 60843;
		16'd13333 : result2 = 61334;
		16'd13334 : result2 = 61844;
		16'd13335 : result2 = 62373;
		16'd13336 : result2 = 62920;
		16'd13337 : result2 = 63484;
		16'd13338 : result2 = 64063;
		16'd13339 : result2 = 64659;
		16'd13340 : result2 = 65269;
		16'd13341 : result2 = 65893;
		16'd13342 : result2 = 66531;
		16'd13343 : result2 = 67182;
		16'd13344 : result2 = 67847;
		16'd13345 : result2 = 68524;
		16'd13346 : result2 = 69214;
		16'd13347 : result2 = 69916;
		16'd13348 : result2 = 70631;
		16'd13349 : result2 = 71357;
		16'd13350 : result2 = 72096;
		16'd13351 : result2 = 72848;
		16'd13352 : result2 = 73611;
		16'd13353 : result2 = 74388;
		16'd13354 : result2 = 75177;
		16'd13355 : result2 = 75979;
		16'd13356 : result2 = 76794;
		16'd13357 : result2 = 77623;
		16'd13358 : result2 = 78466;
		16'd13359 : result2 = 79324;
		16'd13360 : result2 = 80197;
		16'd13361 : result2 = 81086;
		16'd13362 : result2 = 81992;
		16'd13568 : result2 = 55647;
		16'd13569 : result2 = 55278;
		16'd13570 : result2 = 55001;
		16'd13571 : result2 = 54809;
		16'd13572 : result2 = 54692;
		16'd13573 : result2 = 54645;
		16'd13574 : result2 = 54661;
		16'd13575 : result2 = 54734;
		16'd13576 : result2 = 54860;
		16'd13577 : result2 = 55033;
		16'd13578 : result2 = 55250;
		16'd13579 : result2 = 55507;
		16'd13580 : result2 = 55802;
		16'd13581 : result2 = 56130;
		16'd13582 : result2 = 56490;
		16'd13583 : result2 = 56879;
		16'd13584 : result2 = 57295;
		16'd13585 : result2 = 57737;
		16'd13586 : result2 = 58201;
		16'd13587 : result2 = 58688;
		16'd13588 : result2 = 59194;
		16'd13589 : result2 = 59721;
		16'd13590 : result2 = 60265;
		16'd13591 : result2 = 60826;
		16'd13592 : result2 = 61404;
		16'd13593 : result2 = 61997;
		16'd13594 : result2 = 62605;
		16'd13595 : result2 = 63228;
		16'd13596 : result2 = 63863;
		16'd13597 : result2 = 64512;
		16'd13598 : result2 = 65174;
		16'd13599 : result2 = 65849;
		16'd13600 : result2 = 66535;
		16'd13601 : result2 = 67233;
		16'd13602 : result2 = 67944;
		16'd13603 : result2 = 68666;
		16'd13604 : result2 = 69399;
		16'd13605 : result2 = 70144;
		16'd13606 : result2 = 70901;
		16'd13607 : result2 = 71669;
		16'd13608 : result2 = 72449;
		16'd13609 : result2 = 73242;
		16'd13610 : result2 = 74046;
		16'd13611 : result2 = 74863;
		16'd13612 : result2 = 75692;
		16'd13613 : result2 = 76535;
		16'd13614 : result2 = 77392;
		16'd13615 : result2 = 78263;
		16'd13616 : result2 = 79149;
		16'd13617 : result2 = 80051;
		16'd13618 : result2 = 80969;
		16'd13824 : result2 = 52532;
		16'd13825 : result2 = 52301;
		16'd13826 : result2 = 52151;
		16'd13827 : result2 = 52076;
		16'd13828 : result2 = 52067;
		16'd13829 : result2 = 52119;
		16'd13830 : result2 = 52227;
		16'd13831 : result2 = 52386;
		16'd13832 : result2 = 52591;
		16'd13833 : result2 = 52838;
		16'd13834 : result2 = 53124;
		16'd13835 : result2 = 53445;
		16'd13836 : result2 = 53800;
		16'd13837 : result2 = 54185;
		16'd13838 : result2 = 54598;
		16'd13839 : result2 = 55036;
		16'd13840 : result2 = 55499;
		16'd13841 : result2 = 55985;
		16'd13842 : result2 = 56491;
		16'd13843 : result2 = 57017;
		16'd13844 : result2 = 57562;
		16'd13845 : result2 = 58124;
		16'd13846 : result2 = 58702;
		16'd13847 : result2 = 59296;
		16'd13848 : result2 = 59904;
		16'd13849 : result2 = 60527;
		16'd13850 : result2 = 61163;
		16'd13851 : result2 = 61812;
		16'd13852 : result2 = 62474;
		16'd13853 : result2 = 63148;
		16'd13854 : result2 = 63834;
		16'd13855 : result2 = 64531;
		16'd13856 : result2 = 65239;
		16'd13857 : result2 = 65959;
		16'd13858 : result2 = 66689;
		16'd13859 : result2 = 67431;
		16'd13860 : result2 = 68183;
		16'd13861 : result2 = 68946;
		16'd13862 : result2 = 69721;
		16'd13863 : result2 = 70506;
		16'd13864 : result2 = 71303;
		16'd13865 : result2 = 72111;
		16'd13866 : result2 = 72931;
		16'd13867 : result2 = 73762;
		16'd13868 : result2 = 74606;
		16'd13869 : result2 = 75463;
		16'd13870 : result2 = 76334;
		16'd13871 : result2 = 77218;
		16'd13872 : result2 = 78117;
		16'd13873 : result2 = 79031;
		16'd13874 : result2 = 79961;
		16'd14080 : result2 = 49421;
		16'd14081 : result2 = 49331;
		16'd14082 : result2 = 49311;
		16'd14083 : result2 = 49354;
		16'd14084 : result2 = 49455;
		16'd14085 : result2 = 49608;
		16'd14086 : result2 = 49809;
		16'd14087 : result2 = 50053;
		16'd14088 : result2 = 50338;
		16'd14089 : result2 = 50659;
		16'd14090 : result2 = 51014;
		16'd14091 : result2 = 51401;
		16'd14092 : result2 = 51815;
		16'd14093 : result2 = 52257;
		16'd14094 : result2 = 52723;
		16'd14095 : result2 = 53211;
		16'd14096 : result2 = 53721;
		16'd14097 : result2 = 54251;
		16'd14098 : result2 = 54799;
		16'd14099 : result2 = 55365;
		16'd14100 : result2 = 55947;
		16'd14101 : result2 = 56545;
		16'd14102 : result2 = 57157;
		16'd14103 : result2 = 57783;
		16'd14104 : result2 = 58422;
		16'd14105 : result2 = 59074;
		16'd14106 : result2 = 59739;
		16'd14107 : result2 = 60415;
		16'd14108 : result2 = 61102;
		16'd14109 : result2 = 61800;
		16'd14110 : result2 = 62510;
		16'd14111 : result2 = 63230;
		16'd14112 : result2 = 63960;
		16'd14113 : result2 = 64700;
		16'd14114 : result2 = 65451;
		16'd14115 : result2 = 66212;
		16'd14116 : result2 = 66983;
		16'd14117 : result2 = 67765;
		16'd14118 : result2 = 68557;
		16'd14119 : result2 = 69359;
		16'd14120 : result2 = 70172;
		16'd14121 : result2 = 70996;
		16'd14122 : result2 = 71831;
		16'd14123 : result2 = 72678;
		16'd14124 : result2 = 73536;
		16'd14125 : result2 = 74407;
		16'd14126 : result2 = 75291;
		16'd14127 : result2 = 76188;
		16'd14128 : result2 = 77100;
		16'd14129 : result2 = 78026;
		16'd14130 : result2 = 78969;
		16'd14336 : result2 = 46330;
		16'd14337 : result2 = 46382;
		16'd14338 : result2 = 46492;
		16'd14339 : result2 = 46654;
		16'd14340 : result2 = 46864;
		16'd14341 : result2 = 47118;
		16'd14342 : result2 = 47412;
		16'd14343 : result2 = 47743;
		16'd14344 : result2 = 48107;
		16'd14345 : result2 = 48503;
		16'd14346 : result2 = 48927;
		16'd14347 : result2 = 49377;
		16'd14348 : result2 = 49852;
		16'd14349 : result2 = 50350;
		16'd14350 : result2 = 50868;
		16'd14351 : result2 = 51407;
		16'd14352 : result2 = 51964;
		16'd14353 : result2 = 52537;
		16'd14354 : result2 = 53127;
		16'd14355 : result2 = 53733;
		16'd14356 : result2 = 54352;
		16'd14357 : result2 = 54985;
		16'd14358 : result2 = 55631;
		16'd14359 : result2 = 56289;
		16'd14360 : result2 = 56959;
		16'd14361 : result2 = 57640;
		16'd14362 : result2 = 58332;
		16'd14363 : result2 = 59035;
		16'd14364 : result2 = 59748;
		16'd14365 : result2 = 60471;
		16'd14366 : result2 = 61204;
		16'd14367 : result2 = 61946;
		16'd14368 : result2 = 62698;
		16'd14369 : result2 = 63459;
		16'd14370 : result2 = 64230;
		16'd14371 : result2 = 65010;
		16'd14372 : result2 = 65800;
		16'd14373 : result2 = 66600;
		16'd14374 : result2 = 67409;
		16'd14375 : result2 = 68228;
		16'd14376 : result2 = 69057;
		16'd14377 : result2 = 69897;
		16'd14378 : result2 = 70747;
		16'd14379 : result2 = 71609;
		16'd14380 : result2 = 72482;
		16'd14381 : result2 = 73367;
		16'd14382 : result2 = 74264;
		16'd14383 : result2 = 75174;
		16'd14384 : result2 = 76099;
		16'd14385 : result2 = 77038;
		16'd14386 : result2 = 77992;
		16'd14592 : result2 = 43272;
		16'd14593 : result2 = 43465;
		16'd14594 : result2 = 43704;
		16'd14595 : result2 = 43985;
		16'd14596 : result2 = 44304;
		16'd14597 : result2 = 44658;
		16'd14598 : result2 = 45044;
		16'd14599 : result2 = 45460;
		16'd14600 : result2 = 45903;
		16'd14601 : result2 = 46372;
		16'd14602 : result2 = 46865;
		16'd14603 : result2 = 47379;
		16'd14604 : result2 = 47914;
		16'd14605 : result2 = 48467;
		16'd14606 : result2 = 49038;
		16'd14607 : result2 = 49626;
		16'd14608 : result2 = 50229;
		16'd14609 : result2 = 50846;
		16'd14610 : result2 = 51477;
		16'd14611 : result2 = 52122;
		16'd14612 : result2 = 52778;
		16'd14613 : result2 = 53446;
		16'd14614 : result2 = 54126;
		16'd14615 : result2 = 54816;
		16'd14616 : result2 = 55516;
		16'd14617 : result2 = 56226;
		16'd14618 : result2 = 56946;
		16'd14619 : result2 = 57675;
		16'd14620 : result2 = 58413;
		16'd14621 : result2 = 59160;
		16'd14622 : result2 = 59916;
		16'd14623 : result2 = 60681;
		16'd14624 : result2 = 61454;
		16'd14625 : result2 = 62236;
		16'd14626 : result2 = 63027;
		16'd14627 : result2 = 63826;
		16'd14628 : result2 = 64635;
		16'd14629 : result2 = 65452;
		16'd14630 : result2 = 66279;
		16'd14631 : result2 = 67114;
		16'd14632 : result2 = 67960;
		16'd14633 : result2 = 68815;
		16'd14634 : result2 = 69681;
		16'd14635 : result2 = 70557;
		16'd14636 : result2 = 71444;
		16'd14637 : result2 = 72342;
		16'd14638 : result2 = 73253;
		16'd14639 : result2 = 74177;
		16'd14640 : result2 = 75114;
		16'd14641 : result2 = 76065;
		16'd14642 : result2 = 77032;
		16'd14848 : result2 = 40260;
		16'd14849 : result2 = 40593;
		16'd14850 : result2 = 40959;
		16'd14851 : result2 = 41356;
		16'd14852 : result2 = 41781;
		16'd14853 : result2 = 42233;
		16'd14854 : result2 = 42711;
		16'd14855 : result2 = 43210;
		16'd14856 : result2 = 43732;
		16'd14857 : result2 = 44273;
		16'd14858 : result2 = 44833;
		16'd14859 : result2 = 45410;
		16'd14860 : result2 = 46003;
		16'd14861 : result2 = 46612;
		16'd14862 : result2 = 47234;
		16'd14863 : result2 = 47870;
		16'd14864 : result2 = 48519;
		16'd14865 : result2 = 49180;
		16'd14866 : result2 = 49852;
		16'd14867 : result2 = 50534;
		16'd14868 : result2 = 51227;
		16'd14869 : result2 = 51930;
		16'd14870 : result2 = 52642;
		16'd14871 : result2 = 53364;
		16'd14872 : result2 = 54094;
		16'd14873 : result2 = 54833;
		16'd14874 : result2 = 55579;
		16'd14875 : result2 = 56335;
		16'd14876 : result2 = 57098;
		16'd14877 : result2 = 57869;
		16'd14878 : result2 = 58648;
		16'd14879 : result2 = 59435;
		16'd14880 : result2 = 60229;
		16'd14881 : result2 = 61032;
		16'd14882 : result2 = 61842;
		16'd14883 : result2 = 62661;
		16'd14884 : result2 = 63487;
		16'd14885 : result2 = 64322;
		16'd14886 : result2 = 65166;
		16'd14887 : result2 = 66018;
		16'd14888 : result2 = 66879;
		16'd14889 : result2 = 67750;
		16'd14890 : result2 = 68631;
		16'd14891 : result2 = 69521;
		16'd14892 : result2 = 70423;
		16'd14893 : result2 = 71335;
		16'd14894 : result2 = 72259;
		16'd14895 : result2 = 73196;
		16'd14896 : result2 = 74146;
		16'd14897 : result2 = 75109;
		16'd14898 : result2 = 76088;
		16'd15104 : result2 = 37308;
		16'd15105 : result2 = 37775;
		16'd15106 : result2 = 38264;
		16'd15107 : result2 = 38775;
		16'd15108 : result2 = 39304;
		16'd15109 : result2 = 39852;
		16'd15110 : result2 = 40418;
		16'd15111 : result2 = 41000;
		16'd15112 : result2 = 41597;
		16'd15113 : result2 = 42209;
		16'd15114 : result2 = 42835;
		16'd15115 : result2 = 43473;
		16'd15116 : result2 = 44124;
		16'd15117 : result2 = 44786;
		16'd15118 : result2 = 45460;
		16'd15119 : result2 = 46143;
		16'd15120 : result2 = 46837;
		16'd15121 : result2 = 47540;
		16'd15122 : result2 = 48252;
		16'd15123 : result2 = 48972;
		16'd15124 : result2 = 49701;
		16'd15125 : result2 = 50438;
		16'd15126 : result2 = 51183;
		16'd15127 : result2 = 51935;
		16'd15128 : result2 = 52695;
		16'd15129 : result2 = 53461;
		16'd15130 : result2 = 54235;
		16'd15131 : result2 = 55016;
		16'd15132 : result2 = 55804;
		16'd15133 : result2 = 56598;
		16'd15134 : result2 = 57400;
		16'd15135 : result2 = 58208;
		16'd15136 : result2 = 59024;
		16'd15137 : result2 = 59846;
		16'd15138 : result2 = 60676;
		16'd15139 : result2 = 61513;
		16'd15140 : result2 = 62358;
		16'd15141 : result2 = 63211;
		16'd15142 : result2 = 64071;
		16'd15143 : result2 = 64940;
		16'd15144 : result2 = 65817;
		16'd15145 : result2 = 66703;
		16'd15146 : result2 = 67598;
		16'd15147 : result2 = 68503;
		16'd15148 : result2 = 69419;
		16'd15149 : result2 = 70345;
		16'd15150 : result2 = 71282;
		16'd15151 : result2 = 72232;
		16'd15152 : result2 = 73194;
		16'd15153 : result2 = 74170;
		16'd15154 : result2 = 75161;
		16'd15360 : result2 = 34427;
		16'd15361 : result2 = 35023;
		16'd15362 : result2 = 35631;
		16'd15363 : result2 = 36250;
		16'd15364 : result2 = 36880;
		16'd15365 : result2 = 37521;
		16'd15366 : result2 = 38172;
		16'd15367 : result2 = 38833;
		16'd15368 : result2 = 39504;
		16'd15369 : result2 = 40185;
		16'd15370 : result2 = 40874;
		16'd15371 : result2 = 41573;
		16'd15372 : result2 = 42279;
		16'd15373 : result2 = 42994;
		16'd15374 : result2 = 43717;
		16'd15375 : result2 = 44447;
		16'd15376 : result2 = 45184;
		16'd15377 : result2 = 45929;
		16'd15378 : result2 = 46680;
		16'd15379 : result2 = 47437;
		16'd15380 : result2 = 48201;
		16'd15381 : result2 = 48972;
		16'd15382 : result2 = 49748;
		16'd15383 : result2 = 50531;
		16'd15384 : result2 = 51319;
		16'd15385 : result2 = 52113;
		16'd15386 : result2 = 52913;
		16'd15387 : result2 = 53719;
		16'd15388 : result2 = 54531;
		16'd15389 : result2 = 55349;
		16'd15390 : result2 = 56173;
		16'd15391 : result2 = 57003;
		16'd15392 : result2 = 57839;
		16'd15393 : result2 = 58681;
		16'd15394 : result2 = 59530;
		16'd15395 : result2 = 60386;
		16'd15396 : result2 = 61248;
		16'd15397 : result2 = 62118;
		16'd15398 : result2 = 62995;
		16'd15399 : result2 = 63880;
		16'd15400 : result2 = 64772;
		16'd15401 : result2 = 65674;
		16'd15402 : result2 = 66584;
		16'd15403 : result2 = 67503;
		16'd15404 : result2 = 68432;
		16'd15405 : result2 = 69372;
		16'd15406 : result2 = 70322;
		16'd15407 : result2 = 71285;
		16'd15408 : result2 = 72259;
		16'd15409 : result2 = 73248;
		16'd15410 : result2 = 74250;
		16'd15616 : result2 = 31626;
		16'd15617 : result2 = 32346;
		16'd15618 : result2 = 33066;
		16'd15619 : result2 = 33789;
		16'd15620 : result2 = 34515;
		16'd15621 : result2 = 35244;
		16'd15622 : result2 = 35977;
		16'd15623 : result2 = 36715;
		16'd15624 : result2 = 37457;
		16'd15625 : result2 = 38204;
		16'd15626 : result2 = 38955;
		16'd15627 : result2 = 39711;
		16'd15628 : result2 = 40472;
		16'd15629 : result2 = 41238;
		16'd15630 : result2 = 42008;
		16'd15631 : result2 = 42784;
		16'd15632 : result2 = 43564;
		16'd15633 : result2 = 44348;
		16'd15634 : result2 = 45137;
		16'd15635 : result2 = 45931;
		16'd15636 : result2 = 46729;
		16'd15637 : result2 = 47532;
		16'd15638 : result2 = 48340;
		16'd15639 : result2 = 49151;
		16'd15640 : result2 = 49968;
		16'd15641 : result2 = 50789;
		16'd15642 : result2 = 51615;
		16'd15643 : result2 = 52446;
		16'd15644 : result2 = 53281;
		16'd15645 : result2 = 54122;
		16'd15646 : result2 = 54968;
		16'd15647 : result2 = 55818;
		16'd15648 : result2 = 56675;
		16'd15649 : result2 = 57537;
		16'd15650 : result2 = 58404;
		16'd15651 : result2 = 59278;
		16'd15652 : result2 = 60158;
		16'd15653 : result2 = 61045;
		16'd15654 : result2 = 61938;
		16'd15655 : result2 = 62839;
		16'd15656 : result2 = 63747;
		16'd15657 : result2 = 64663;
		16'd15658 : result2 = 65587;
		16'd15659 : result2 = 66521;
		16'd15660 : result2 = 67464;
		16'd15661 : result2 = 68417;
		16'd15662 : result2 = 69380;
		16'd15663 : result2 = 70355;
		16'd15664 : result2 = 71342;
		16'd15665 : result2 = 72343;
		16'd15666 : result2 = 73357;
		16'd15872 : result2 = 28916;
		16'd15873 : result2 = 29751;
		16'd15874 : result2 = 30577;
		16'd15875 : result2 = 31398;
		16'd15876 : result2 = 32214;
		16'd15877 : result2 = 33028;
		16'd15878 : result2 = 33839;
		16'd15879 : result2 = 34649;
		16'd15880 : result2 = 35459;
		16'd15881 : result2 = 36269;
		16'd15882 : result2 = 37080;
		16'd15883 : result2 = 37892;
		16'd15884 : result2 = 38705;
		16'd15885 : result2 = 39520;
		16'd15886 : result2 = 40336;
		16'd15887 : result2 = 41155;
		16'd15888 : result2 = 41976;
		16'd15889 : result2 = 42800;
		16'd15890 : result2 = 43626;
		16'd15891 : result2 = 44455;
		16'd15892 : result2 = 45286;
		16'd15893 : result2 = 46121;
		16'd15894 : result2 = 46958;
		16'd15895 : result2 = 47799;
		16'd15896 : result2 = 48643;
		16'd15897 : result2 = 49491;
		16'd15898 : result2 = 50342;
		16'd15899 : result2 = 51196;
		16'd15900 : result2 = 52055;
		16'd15901 : result2 = 52918;
		16'd15902 : result2 = 53785;
		16'd15903 : result2 = 54656;
		16'd15904 : result2 = 55532;
		16'd15905 : result2 = 56413;
		16'd15906 : result2 = 57299;
		16'd15907 : result2 = 58191;
		16'd15908 : result2 = 59088;
		16'd15909 : result2 = 59991;
		16'd15910 : result2 = 60901;
		16'd15911 : result2 = 61817;
		16'd15912 : result2 = 62740;
		16'd15913 : result2 = 63671;
		16'd15914 : result2 = 64610;
		16'd15915 : result2 = 65557;
		16'd15916 : result2 = 66513;
		16'd15917 : result2 = 67479;
		16'd15918 : result2 = 68456;
		16'd15919 : result2 = 69443;
		16'd15920 : result2 = 70443;
		16'd15921 : result2 = 71455;
		16'd15922 : result2 = 72482;
		16'd16128 : result2 = 26304;
		16'd16129 : result2 = 27245;
		16'd16130 : result2 = 28170;
		16'd16131 : result2 = 29082;
		16'd16132 : result2 = 29984;
		16'd16133 : result2 = 30876;
		16'd16134 : result2 = 31761;
		16'd16135 : result2 = 32640;
		16'd16136 : result2 = 33515;
		16'd16137 : result2 = 34385;
		16'd16138 : result2 = 35252;
		16'd16139 : result2 = 36117;
		16'd16140 : result2 = 36980;
		16'd16141 : result2 = 37842;
		16'd16142 : result2 = 38703;
		16'd16143 : result2 = 39564;
		16'd16144 : result2 = 40424;
		16'd16145 : result2 = 41286;
		16'd16146 : result2 = 42147;
		16'd16147 : result2 = 43010;
		16'd16148 : result2 = 43874;
		16'd16149 : result2 = 44739;
		16'd16150 : result2 = 45606;
		16'd16151 : result2 = 46474;
		16'd16152 : result2 = 47345;
		16'd16153 : result2 = 48218;
		16'd16154 : result2 = 49094;
		16'd16155 : result2 = 49972;
		16'd16156 : result2 = 50853;
		16'd16157 : result2 = 51737;
		16'd16158 : result2 = 52625;
		16'd16159 : result2 = 53517;
		16'd16160 : result2 = 54412;
		16'd16161 : result2 = 55312;
		16'd16162 : result2 = 56216;
		16'd16163 : result2 = 57125;
		16'd16164 : result2 = 58039;
		16'd16165 : result2 = 58958;
		16'd16166 : result2 = 59883;
		16'd16167 : result2 = 60815;
		16'd16168 : result2 = 61753;
		16'd16169 : result2 = 62698;
		16'd16170 : result2 = 63651;
		16'd16171 : result2 = 64612;
		16'd16172 : result2 = 65582;
		16'd16173 : result2 = 66561;
		16'd16174 : result2 = 67550;
		16'd16175 : result2 = 68550;
		16'd16176 : result2 = 69561;
		16'd16177 : result2 = 70586;
		16'd16178 : result2 = 71624;
		16'd16384 : result2 = 23795;
		16'd16385 : result2 = 24833;
		16'd16386 : result2 = 25850;
		16'd16387 : result2 = 26847;
		16'd16388 : result2 = 27827;
		16'd16389 : result2 = 28793;
		16'd16390 : result2 = 29747;
		16'd16391 : result2 = 30691;
		16'd16392 : result2 = 31626;
		16'd16393 : result2 = 32553;
		16'd16394 : result2 = 33474;
		16'd16395 : result2 = 34389;
		16'd16396 : result2 = 35300;
		16'd16397 : result2 = 36206;
		16'd16398 : result2 = 37110;
		16'd16399 : result2 = 38011;
		16'd16400 : result2 = 38909;
		16'd16401 : result2 = 39807;
		16'd16402 : result2 = 40703;
		16'd16403 : result2 = 41598;
		16'd16404 : result2 = 42493;
		16'd16405 : result2 = 43387;
		16'd16406 : result2 = 44283;
		16'd16407 : result2 = 45178;
		16'd16408 : result2 = 46075;
		16'd16409 : result2 = 46973;
		16'd16410 : result2 = 47872;
		16'd16411 : result2 = 48773;
		16'd16412 : result2 = 49676;
		16'd16413 : result2 = 50581;
		16'd16414 : result2 = 51489;
		16'd16415 : result2 = 52400;
		16'd16416 : result2 = 53315;
		16'd16417 : result2 = 54232;
		16'd16418 : result2 = 55154;
		16'd16419 : result2 = 56080;
		16'd16420 : result2 = 57010;
		16'd16421 : result2 = 57946;
		16'd16422 : result2 = 58886;
		16'd16423 : result2 = 59833;
		16'd16424 : result2 = 60785;
		16'd16425 : result2 = 61745;
		16'd16426 : result2 = 62712;
		16'd16427 : result2 = 63686;
		16'd16428 : result2 = 64669;
		16'd16429 : result2 = 65661;
		16'd16430 : result2 = 66662;
		16'd16431 : result2 = 67675;
		16'd16432 : result2 = 68698;
		16'd16433 : result2 = 69735;
		16'd16434 : result2 = 70784;
		16'd16640 : result2 = 21393;
		16'd16641 : result2 = 22520;
		16'd16642 : result2 = 23620;
		16'd16643 : result2 = 24694;
		16'd16644 : result2 = 25748;
		16'd16645 : result2 = 26782;
		16'd16646 : result2 = 27800;
		16'd16647 : result2 = 28804;
		16'd16648 : result2 = 29796;
		16'd16649 : result2 = 30777;
		16'd16650 : result2 = 31748;
		16'd16651 : result2 = 32710;
		16'd16652 : result2 = 33666;
		16'd16653 : result2 = 34615;
		16'd16654 : result2 = 35559;
		16'd16655 : result2 = 36498;
		16'd16656 : result2 = 37433;
		16'd16657 : result2 = 38365;
		16'd16658 : result2 = 39293;
		16'd16659 : result2 = 40220;
		16'd16660 : result2 = 41144;
		16'd16661 : result2 = 42068;
		16'd16662 : result2 = 42990;
		16'd16663 : result2 = 43912;
		16'd16664 : result2 = 44833;
		16'd16665 : result2 = 45755;
		16'd16666 : result2 = 46677;
		16'd16667 : result2 = 47600;
		16'd16668 : result2 = 48524;
		16'd16669 : result2 = 49450;
		16'd16670 : result2 = 50378;
		16'd16671 : result2 = 51308;
		16'd16672 : result2 = 52240;
		16'd16673 : result2 = 53176;
		16'd16674 : result2 = 54115;
		16'd16675 : result2 = 55057;
		16'd16676 : result2 = 56003;
		16'd16677 : result2 = 56954;
		16'd16678 : result2 = 57910;
		16'd16679 : result2 = 58871;
		16'd16680 : result2 = 59838;
		16'd16681 : result2 = 60812;
		16'd16682 : result2 = 61792;
		16'd16683 : result2 = 62779;
		16'd16684 : result2 = 63775;
		16'd16685 : result2 = 64780;
		16'd16686 : result2 = 65794;
		16'd16687 : result2 = 66818;
		16'd16688 : result2 = 67854;
		16'd16689 : result2 = 68901;
		16'd16690 : result2 = 69963;
		16'd16896 : result2 = 19102;
		16'd16897 : result2 = 20309;
		16'd16898 : result2 = 21483;
		16'd16899 : result2 = 22628;
		16'd16900 : result2 = 23748;
		16'd16901 : result2 = 24845;
		16'd16902 : result2 = 25922;
		16'd16903 : result2 = 26982;
		16'd16904 : result2 = 28026;
		16'd16905 : result2 = 29057;
		16'd16906 : result2 = 30075;
		16'd16907 : result2 = 31082;
		16'd16908 : result2 = 32080;
		16'd16909 : result2 = 33069;
		16'd16910 : result2 = 34051;
		16'd16911 : result2 = 35027;
		16'd16912 : result2 = 35996;
		16'd16913 : result2 = 36960;
		16'd16914 : result2 = 37921;
		16'd16915 : result2 = 38877;
		16'd16916 : result2 = 39830;
		16'd16917 : result2 = 40781;
		16'd16918 : result2 = 41729;
		16'd16919 : result2 = 42676;
		16'd16920 : result2 = 43621;
		16'd16921 : result2 = 44566;
		16'd16922 : result2 = 45510;
		16'd16923 : result2 = 46455;
		16'd16924 : result2 = 47399;
		16'd16925 : result2 = 48345;
		16'd16926 : result2 = 49292;
		16'd16927 : result2 = 50240;
		16'd16928 : result2 = 51190;
		16'd16929 : result2 = 52143;
		16'd16930 : result2 = 53098;
		16'd16931 : result2 = 54057;
		16'd16932 : result2 = 55019;
		16'd16933 : result2 = 55985;
		16'd16934 : result2 = 56955;
		16'd16935 : result2 = 57931;
		16'd16936 : result2 = 58912;
		16'd16937 : result2 = 59899;
		16'd16938 : result2 = 60892;
		16'd16939 : result2 = 61893;
		16'd16940 : result2 = 62901;
		16'd16941 : result2 = 63918;
		16'd16942 : result2 = 64944;
		16'd16943 : result2 = 65980;
		16'd16944 : result2 = 67027;
		16'd16945 : result2 = 68087;
		16'd16946 : result2 = 69159;
		16'd17152 : result2 = 16923;
		16'd17153 : result2 = 18200;
		16'd17154 : result2 = 19441;
		16'd17155 : result2 = 20650;
		16'd17156 : result2 = 21830;
		16'd17157 : result2 = 22984;
		16'd17158 : result2 = 24115;
		16'd17159 : result2 = 25226;
		16'd17160 : result2 = 26319;
		16'd17161 : result2 = 27396;
		16'd17162 : result2 = 28457;
		16'd17163 : result2 = 29506;
		16'd17164 : result2 = 30544;
		16'd17165 : result2 = 31571;
		16'd17166 : result2 = 32588;
		16'd17167 : result2 = 33598;
		16'd17168 : result2 = 34600;
		16'd17169 : result2 = 35595;
		16'd17170 : result2 = 36585;
		16'd17171 : result2 = 37570;
		16'd17172 : result2 = 38550;
		16'd17173 : result2 = 39527;
		16'd17174 : result2 = 40500;
		16'd17175 : result2 = 41471;
		16'd17176 : result2 = 42439;
		16'd17177 : result2 = 43406;
		16'd17178 : result2 = 44372;
		16'd17179 : result2 = 45336;
		16'd17180 : result2 = 46301;
		16'd17181 : result2 = 47266;
		16'd17182 : result2 = 48231;
		16'd17183 : result2 = 49197;
		16'd17184 : result2 = 50164;
		16'd17185 : result2 = 51134;
		16'd17186 : result2 = 52105;
		16'd17187 : result2 = 53079;
		16'd17188 : result2 = 54056;
		16'd17189 : result2 = 55037;
		16'd17190 : result2 = 56022;
		16'd17191 : result2 = 57012;
		16'd17192 : result2 = 58006;
		16'd17193 : result2 = 59006;
		16'd17194 : result2 = 60013;
		16'd17195 : result2 = 61026;
		16'd17196 : result2 = 62047;
		16'd17197 : result2 = 63076;
		16'd17198 : result2 = 64114;
		16'd17199 : result2 = 65162;
		16'd17200 : result2 = 66220;
		16'd17201 : result2 = 67291;
		16'd17202 : result2 = 68374;
		16'd17408 : result2 = 14856;
		16'd17409 : result2 = 16195;
		16'd17410 : result2 = 17495;
		16'd17411 : result2 = 18760;
		16'd17412 : result2 = 19994;
		16'd17413 : result2 = 21200;
		16'd17414 : result2 = 22380;
		16'd17415 : result2 = 23538;
		16'd17416 : result2 = 24675;
		16'd17417 : result2 = 25794;
		16'd17418 : result2 = 26896;
		16'd17419 : result2 = 27984;
		16'd17420 : result2 = 29058;
		16'd17421 : result2 = 30120;
		16'd17422 : result2 = 31171;
		16'd17423 : result2 = 32213;
		16'd17424 : result2 = 33245;
		16'd17425 : result2 = 34270;
		16'd17426 : result2 = 35288;
		16'd17427 : result2 = 36300;
		16'd17428 : result2 = 37306;
		16'd17429 : result2 = 38307;
		16'd17430 : result2 = 39304;
		16'd17431 : result2 = 40298;
		16'd17432 : result2 = 41288;
		16'd17433 : result2 = 42276;
		16'd17434 : result2 = 43262;
		16'd17435 : result2 = 44246;
		16'd17436 : result2 = 45230;
		16'd17437 : result2 = 46213;
		16'd17438 : result2 = 47196;
		16'd17439 : result2 = 48179;
		16'd17440 : result2 = 49163;
		16'd17441 : result2 = 50148;
		16'd17442 : result2 = 51136;
		16'd17443 : result2 = 52125;
		16'd17444 : result2 = 53117;
		16'd17445 : result2 = 54112;
		16'd17446 : result2 = 55111;
		16'd17447 : result2 = 56114;
		16'd17448 : result2 = 57122;
		16'd17449 : result2 = 58135;
		16'd17450 : result2 = 59154;
		16'd17451 : result2 = 60180;
		16'd17452 : result2 = 61212;
		16'd17453 : result2 = 62253;
		16'd17454 : result2 = 63303;
		16'd17455 : result2 = 64362;
		16'd17456 : result2 = 65432;
		16'd17457 : result2 = 66514;
		16'd17458 : result2 = 67607;
		16'd17664 : result2 = 12901;
		16'd17665 : result2 = 14294;
		16'd17666 : result2 = 15645;
		16'd17667 : result2 = 16960;
		16'd17668 : result2 = 18242;
		16'd17669 : result2 = 19493;
		16'd17670 : result2 = 20718;
		16'd17671 : result2 = 21918;
		16'd17672 : result2 = 23095;
		16'd17673 : result2 = 24253;
		16'd17674 : result2 = 25393;
		16'd17675 : result2 = 26516;
		16'd17676 : result2 = 27624;
		16'd17677 : result2 = 28718;
		16'd17678 : result2 = 29801;
		16'd17679 : result2 = 30872;
		16'd17680 : result2 = 31933;
		16'd17681 : result2 = 32986;
		16'd17682 : result2 = 34030;
		16'd17683 : result2 = 35067;
		16'd17684 : result2 = 36097;
		16'd17685 : result2 = 37122;
		16'd17686 : result2 = 38142;
		16'd17687 : result2 = 39157;
		16'd17688 : result2 = 40168;
		16'd17689 : result2 = 41176;
		16'd17690 : result2 = 42182;
		16'd17691 : result2 = 43185;
		16'd17692 : result2 = 44187;
		16'd17693 : result2 = 45187;
		16'd17694 : result2 = 46187;
		16'd17695 : result2 = 47187;
		16'd17696 : result2 = 48187;
		16'd17697 : result2 = 49188;
		16'd17698 : result2 = 50190;
		16'd17699 : result2 = 51194;
		16'd17700 : result2 = 52200;
		16'd17701 : result2 = 53210;
		16'd17702 : result2 = 54222;
		16'd17703 : result2 = 55238;
		16'd17704 : result2 = 56259;
		16'd17705 : result2 = 57285;
		16'd17706 : result2 = 58316;
		16'd17707 : result2 = 59354;
		16'd17708 : result2 = 60398;
		16'd17709 : result2 = 61451;
		16'd17710 : result2 = 62512;
		16'd17711 : result2 = 63582;
		16'd17712 : result2 = 64663;
		16'd17713 : result2 = 65755;
		16'd17714 : result2 = 66859;
		16'd17920 : result2 = 11056;
		16'd17921 : result2 = 12494;
		16'd17922 : result2 = 13890;
		16'd17923 : result2 = 15249;
		16'd17924 : result2 = 16572;
		16'd17925 : result2 = 17864;
		16'd17926 : result2 = 19128;
		16'd17927 : result2 = 20366;
		16'd17928 : result2 = 21580;
		16'd17929 : result2 = 22773;
		16'd17930 : result2 = 23947;
		16'd17931 : result2 = 25102;
		16'd17932 : result2 = 26241;
		16'd17933 : result2 = 27366;
		16'd17934 : result2 = 28477;
		16'd17935 : result2 = 29576;
		16'd17936 : result2 = 30664;
		16'd17937 : result2 = 31742;
		16'd17938 : result2 = 32811;
		16'd17939 : result2 = 33872;
		16'd17940 : result2 = 34926;
		16'd17941 : result2 = 35972;
		16'd17942 : result2 = 37013;
		16'd17943 : result2 = 38049;
		16'd17944 : result2 = 39080;
		16'd17945 : result2 = 40108;
		16'd17946 : result2 = 41132;
		16'd17947 : result2 = 42153;
		16'd17948 : result2 = 43172;
		16'd17949 : result2 = 44189;
		16'd17950 : result2 = 45206;
		16'd17951 : result2 = 46221;
		16'd17952 : result2 = 47237;
		16'd17953 : result2 = 48252;
		16'd17954 : result2 = 49269;
		16'd17955 : result2 = 50287;
		16'd17956 : result2 = 51307;
		16'd17957 : result2 = 52330;
		16'd17958 : result2 = 53356;
		16'd17959 : result2 = 54385;
		16'd17960 : result2 = 55418;
		16'd17961 : result2 = 56456;
		16'd17962 : result2 = 57499;
		16'd17963 : result2 = 58549;
		16'd17964 : result2 = 59605;
		16'd17965 : result2 = 60669;
		16'd17966 : result2 = 61741;
		16'd17967 : result2 = 62822;
		16'd17968 : result2 = 63913;
		16'd17969 : result2 = 65015;
		16'd17970 : result2 = 66127;

    16'd19758 : result2 = 55500;
endcase;
end

endmodule
